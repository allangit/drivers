
.subckt AND2X1 IN1 IN2 Q VDD VSS
mmp2 net1 IN2 VDD VDD p12 l = 0.1u w = 0.41u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.41u m = 1
mmp3 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 Q net1 VSS VSS n12 l = 0.1u w = 0.4u m = 1


.ends AND2X1



.subckt AND2X2 IN1 IN2 Q VDD VSS
mmp4 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp5 net1 IN1 VDD VDD p12 l = 0.1u w = 0.41u m = 1
mmp6 net1 IN2 VDD VDD p12 l = 0.1u w = 0.41u m = 1
mmn4 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net1 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 Q net1 VSS VSS n12 l = 0.1u w = 0.4u m = 2


.ends AND2X2



.subckt AND2X4 IN1 IN2 Q VDD VSS
mmp4 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmp5 net1 IN1 VDD VDD p12 l = 0.1u w = 0.41u m = 1
mmp6 net1 IN2 VDD VDD p12 l = 0.1u w = 0.41u m = 1
mmn4 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net1 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 Q net1 VSS VSS n12 l = 0.1u w = 0.4u m = 4


.ends AND2X4



.subckt AND3X1 IN1 IN2 IN3 Q VDD VSS
mmn2 net2 IN2 net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net3 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 Q net1 VSS VSS n12 l = 0.1u w = 0.38u m = 1
mmp2 net1 IN2 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp3 net1 IN3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp4 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 1


.ends AND3X1



.subckt AND3X2 IN1 IN2 IN3 Q VDD VSS
mmn5 net2 IN2 net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net3 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net1 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 Q net1 VSS VSS n12 l = 0.1u w = 0.36u m = 2
mmp5 net1 IN3 VDD VDD p12 l = 0.1u w = 0.31u m = 1
mmp6 net1 IN1 VDD VDD p12 l = 0.1u w = 0.31u m = 1
mmp7 net1 IN2 VDD VDD p12 l = 0.1u w = 0.31u m = 1
mmp8 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 2


.ends AND3X2



.subckt AND3X4 IN1 IN2 IN3 Q VDD VSS
mmn5 net2 IN2 net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net3 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net1 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 Q net1 VSS VSS n12 l = 0.1u w = 0.36u m = 4
mmp5 net1 IN3 VDD VDD p12 l = 0.1u w = 0.31u m = 1
mmp6 net1 IN1 VDD VDD p12 l = 0.1u w = 0.31u m = 1
mmp7 net1 IN2 VDD VDD p12 l = 0.1u w = 0.31u m = 1
mmp8 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 4


.ends AND3X4



.subckt AND4X1 IN1 IN2 IN3 IN4 Q VDD VSS
mmn2 net2 IN2 net3 VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 net3 IN3 net4 VSS n12 l = 0.1u w = 0.24u m = 1
mmn1 net1 IN1 net2 VSS n12 l = 0.1u w = 0.24u m = 1
mmn4 net4 IN4 VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn5 Q net1 VSS VSS n12 l = 0.1u w = 0.35u m = 1
mmp2 net1 IN2 VDD VDD p12 l = 0.1u w = 0.28u m = 1
mmp3 net1 IN3 VDD VDD p12 l = 0.1u w = 0.28u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.28u m = 1
mmp4 net1 IN4 VDD VDD p12 l = 0.1u w = 0.28u m = 1
mmp5 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 1


.ends AND4X1



.subckt AND4X2 IN1 IN2 IN3 IN4 Q VDD VSS
mmp6 net1 IN3 VDD VDD p12 l = 0.1u w = 0.28u m = 1
mmp7 net1 IN1 VDD VDD p12 l = 0.1u w = 0.28u m = 1
mmp8 net1 IN4 VDD VDD p12 l = 0.1u w = 0.28u m = 1
mmp9 net1 IN2 VDD VDD p12 l = 0.1u w = 0.28u m = 1
mmp10 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmn6 net2 IN2 net3 VSS n12 l = 0.1u w = 0.26u m = 1
mmn7 net3 IN3 net4 VSS n12 l = 0.1u w = 0.26u m = 1
mmn8 net1 IN1 net2 VSS n12 l = 0.1u w = 0.26u m = 1
mmn9 net4 IN4 VSS VSS n12 l = 0.1u w = 0.26u m = 1
mmn10 Q net1 VSS VSS n12 l = 0.1u w = 0.38u m = 2


.ends AND4X2



.subckt AND4X4 IN1 IN2 IN3 IN4 Q VDD VSS
mmp6 net1 IN3 VDD VDD p12 l = 0.1u w = 0.28u m = 1
mmp7 net1 IN1 VDD VDD p12 l = 0.1u w = 0.28u m = 1
mmp8 net1 IN4 VDD VDD p12 l = 0.1u w = 0.28u m = 1
mmp9 net1 IN2 VDD VDD p12 l = 0.1u w = 0.28u m = 1
mmp10 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmn6 net2 IN2 net3 VSS n12 l = 0.1u w = 0.26u m = 1
mmn7 net3 IN3 net4 VSS n12 l = 0.1u w = 0.26u m = 1
mmn8 net1 IN1 net2 VSS n12 l = 0.1u w = 0.26u m = 1
mmn9 net4 IN4 VSS VSS n12 l = 0.1u w = 0.26u m = 1
mmn10 Q net1 VSS VSS n12 l = 0.1u w = 0.42u m = 4


.ends AND4X4



.subckt ANTENNA INP VDD VSS





.ends ANTENNA




.subckt AO21X1 IN1 IN2 IN3 Q VDD VSS
mmp4 Q net3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.54u m = 1
mmp3 net3 IN3 net1 VDD p12 l = 0.1u w = 0.65u m = 1
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.54u m = 1
mmn2 net3 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net3 IN3 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn4 Q net3 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends AO21X1



.subckt AO21X2 IN1 IN2 IN3 Q VDD VSS
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net3 IN3 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn4 Q net3 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn2 net3 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.54u m = 1
mmp4 Q net3 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.54u m = 1
mmp3 net3 IN3 net1 VDD p12 l = 0.1u w = 0.65u m = 1


.ends AO21X2



.subckt AO221X1 IN1 IN2 IN3 IN4 IN5 Q VDD VSS
mmn4 net5 IN3 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 Q net5 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn3 net4 IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 IN5 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn2 net5 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmp3 net3 IN4 net1 VDD p12 l = 0.1u w = 0.58u m = 1
mmp6 Q net5 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp4 net3 IN3 net1 VDD p12 l = 0.1u w = 0.58u m = 1
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.58u m = 1
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.58u m = 1
mmp5 net5 IN5 net3 VDD p12 l = 0.1u w = 0.9u m = 1


.ends AO221X1



.subckt AO221X2 IN1 IN2 IN3 IN4 IN5 Q VDD VSS
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.58u m = 1
mmp3 net3 IN4 net1 VDD p12 l = 0.1u w = 0.58u m = 1
mmp5 net5 IN5 net3 VDD p12 l = 0.1u w = 0.9u m = 1
mmp6 Q net5 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.58u m = 1
mmp4 net3 IN3 net1 VDD p12 l = 0.1u w = 0.58u m = 1
mmn4 net5 IN3 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 Q net5 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 IN5 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn2 net5 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net4 IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends AO221X2



.subckt AO222X1 IN1 IN2 IN3 IN4 IN5 IN6 Q VDD VSS
mmp5 net5 IN6 net3 VDD p12 l = 0.1u w = 0.62u m = 1
mmp4 net3 IN3 net1 VDD p12 l = 0.1u w = 0.62u m = 1
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp3 net3 IN4 net1 VDD p12 l = 0.1u w = 0.62u m = 1
mmp6 net5 IN5 net3 VDD p12 l = 0.1u w = 0.62u m = 1
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp7 Q net5 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net5 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net5 IN5 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net4 IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net5 IN3 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net6 IN6 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 Q net5 VSS VSS n12 l = 0.1u w = 0.43u m = 1


.ends AO222X1



.subckt AO222X2 IN1 IN2 IN3 IN4 IN5 IN6 Q VDD VSS
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp5 net5 IN6 net3 VDD p12 l = 0.1u w = 0.62u m = 1
mmp3 net3 IN4 net1 VDD p12 l = 0.1u w = 0.62u m = 1
mmp4 net3 IN3 net1 VDD p12 l = 0.1u w = 0.62u m = 1
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp7 Q net5 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp6 net5 IN5 net3 VDD p12 l = 0.1u w = 0.62u m = 1
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net5 IN5 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 Q net5 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn4 net5 IN3 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net6 IN6 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net5 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net4 IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends AO222X2



.subckt AO22X1 IN1 IN2 IN3 IN4 Q VDD VSS
mmn2 net3 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net3 IN3 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 Q net3 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn3 net4 IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp3 net3 IN4 net1 VDD p12 l = 0.1u w = 0.47u m = 1
mmp5 Q net3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.47u m = 1
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.47u m = 1
mmp4 net3 IN3 net1 VDD p12 l = 0.1u w = 0.47u m = 1


.ends AO22X1



.subckt AO22X2 IN1 IN2 IN3 IN4 Q VDD VSS
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.47u m = 1
mmp5 Q net3 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.47u m = 1
mmp3 net3 IN4 net1 VDD p12 l = 0.1u w = 0.47u m = 1
mmp4 net3 IN3 net1 VDD p12 l = 0.1u w = 0.47u m = 1
mmn2 net3 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net4 IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net3 IN3 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 Q net3 VSS VSS n12 l = 0.1u w = 0.43u m = 2


.ends AO22X2



.subckt AOBUFX1 INP VDD VDDG VSS Z
mmn2 Z netp1 VSS VSS n12 l = 0.1u w = 0.49u m = 1
mmn1 netp1 INP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 Z netp1 VDDG VDDG p12 l = 0.1u w = 1.12u m = 1
mmp1 netp1 INP VDDG VDDG p12 l = 0.1u w = 0.5u m = 1


.ends AOBUFX1



.subckt AOBUFX2 INP VDD VDDG VSS Z
mmn2 Z netp1 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn1 netp1 INP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 Z netp1 VDDG VDDG p12 l = 0.1u w = 2.2u m = 1
mmp1 netp1 INP VDDG VDDG p12 l = 0.1u w = 0.55u m = 1


.ends AOBUFX2



.subckt AOBUFX4 INP VDD VDDG VSS Z
mmn2 Z netp1 VSS VSS n12 l = 0.1u w = 1.9u m = 1
mmn1 netp1 INP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 Z netp1 VDDG VDDG p12 l = 0.1u w = 4.2u m = 1
mmp1 netp1 INP VDDG VDDG p12 l = 0.1u w = 0.6u m = 1


.ends AOBUFX4



.subckt AODFFARX1 CLK D Q QN RSTB VDD VDDG VSS
mmp03 net06 D VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDDG VDDG p12 l = 0.1u w = 1.12u m = 1
mmp12 net7 net8 net10 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDDG VDDG p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKP VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP net06 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDDG VDDG p12 l = 0.1u w = 1.12u m = 1
mmp7 net7 CLKN net2 VDDG p12 l = 0.1u w = 0.45u m = 1
mmp8 net8 net7 VDDG VDDG p12 l = 0.1u w = 0.39u m = 1
mmp6 net1 net2 net4 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDDG VDDG p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDDG VDDG p12 l = 0.1u w = 0.39u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.44u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends AODFFARX1



.subckt AODFFARX2 CLK D Q QN RSTB VDD VDDG VSS
mmp03 net06 D VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDDG VDDG p12 l = 0.1u w = 2.2u m = 1
mmp12 net7 net8 net10 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDDG VDDG p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKP VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP net06 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDDG VDDG p12 l = 0.1u w = 2.24u m = 1
mmp7 net7 CLKN net2 VDDG p12 l = 0.1u w = 0.45u m = 1
mmp8 net8 net7 VDDG VDDG p12 l = 0.1u w = 0.39u m = 1
mmp6 net1 net2 net4 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDDG VDDG p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDDG VDDG p12 l = 0.1u w = 0.39u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.76u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends AODFFARX2



.subckt AODFFNARX1 CLK D Q QN RSTB VDD VDDG VSS
mmp03 net06 D VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDDG VDDG p12 l = 0.1u w = 1.1u m = 1
mmp12 net7 net8 net10 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDDG VDDG p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKN VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKN net06 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDDG VDDG p12 l = 0.1u w = 1.12u m = 1
mmp7 net7 CLKP net2 VDDG p12 l = 0.1u w = 0.62u m = 1
mmp8 net8 net7 VDDG VDDG p12 l = 0.1u w = 0.39u m = 1
mmp6 net1 net2 net4 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDDG VDDG p12 l = 0.1u w = 0.44u m = 1
mmp9 net8 RSTB VDDG VDDG p12 l = 0.1u w = 0.39u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.44u m = 1


.ends AODFFNARX1



.subckt AODFFNARX2 CLK D Q QN RSTB VDD VDDG VSS
mmp03 net06 D VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDDG VDDG p12 l = 0.1u w = 1u m = 2
mmp12 net7 net8 net10 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDDG VDDG p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKN VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKN net06 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDDG VDDG p12 l = 0.1u w = 1.12u m = 2
mmp7 net7 CLKP net2 VDDG p12 l = 0.1u w = 0.62u m = 1
mmp8 net8 net7 VDDG VDDG p12 l = 0.1u w = 0.39u m = 1
mmp6 net1 net2 net4 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDDG p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDDG VDDG p12 l = 0.1u w = 0.44u m = 1
mmp9 net8 RSTB VDDG VDDG p12 l = 0.1u w = 0.39u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.44u m = 2
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.56u m = 2
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.44u m = 1


.ends AODFFNARX2



.subckt AOI21X1 IN1 IN2 IN3 QN VDD VSS
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp3 net3 IN3 net1 VDD p12 l = 0.1u w = 0.65u m = 1
mmp5 QN net4 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp4 net4 net3 VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmn5 QN net4 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn3 net3 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net4 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends AOI21X1



.subckt AOI21X2 IN1 IN2 IN3 QN VDD VSS
mmp3 net3 IN3 net1 VDD p12 l = 0.1u w = 0.65u m = 1
mmp4 net4 net3 VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp5 QN net4 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmn2 net3 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net4 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 QN net4 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn3 net3 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends AOI21X2



.subckt AOI221X1 IN1 IN2 IN3 IN4 IN5 QN VDD VSS
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net4 IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 IN5 VSS VSS n12 l = 0.1u w = 0.17u m = 1
mmn4 net5 IN3 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net5 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net6 net5 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 QN net6 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmp5 net5 IN5 net3 VDD p12 l = 0.1u w = 0.99u m = 1
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp4 net3 IN3 net1 VDD p12 l = 0.1u w = 0.47u m = 1
mmp3 net3 IN4 net1 VDD p12 l = 0.1u w = 0.47u m = 1
mmp7 QN net6 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp6 net6 net5 VDD VDD p12 l = 0.1u w = 0.5u m = 1


.ends AOI221X1



.subckt AOI221X2 IN1 IN2 IN3 IN4 IN5 QN VDD VSS
mmn6 net6 net5 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 QN net6 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn5 net5 IN5 VSS VSS n12 l = 0.1u w = 0.17u m = 1
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net5 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net4 IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net5 IN3 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp5 net5 IN5 net3 VDD p12 l = 0.1u w = 0.99u m = 1
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp6 net6 net5 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp3 net3 IN4 net1 VDD p12 l = 0.1u w = 0.47u m = 1
mmp4 net3 IN3 net1 VDD p12 l = 0.1u w = 0.47u m = 1
mmp7 QN net6 VDD VDD p12 l = 0.1u w = 1.12u m = 2


.ends AOI221X2



.subckt AOI222X1 IN1 IN2 IN3 IN4 IN5 IN6 QN VDD VSS
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp4 net3 IN3 net1 VDD p12 l = 0.1u w = 0.55u m = 1
mmp6 net6 IN5 net3 VDD p12 l = 0.1u w = 0.55u m = 1
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp3 net3 IN4 net1 VDD p12 l = 0.1u w = 0.55u m = 1
mmp5 net6 IN6 net3 VDD p12 l = 0.1u w = 0.55u m = 1
mmp7 net7 net6 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp8 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net4 IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 IN6 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net6 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 IN3 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net6 IN5 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 net6 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 QN net7 VSS VSS n12 l = 0.1u w = 0.43u m = 1


.ends AOI222X1



.subckt AOI222X2 IN1 IN2 IN3 IN4 IN5 IN6 QN VDD VSS
mmn2 net6 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 net6 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net4 IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 IN3 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 IN6 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net6 IN5 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 QN net7 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmp5 net6 IN6 net3 VDD p12 l = 0.1u w = 0.55u m = 1
mmp3 net3 IN4 net1 VDD p12 l = 0.1u w = 0.55u m = 1
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp6 net6 IN5 net3 VDD p12 l = 0.1u w = 0.55u m = 1
mmp8 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp7 net7 net6 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp4 net3 IN3 net1 VDD p12 l = 0.1u w = 0.55u m = 1


.ends AOI222X2



.subckt AOI22X1 IN1 IN2 IN3 IN4 QN VDD VSS
mmp5 net5 net3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp4 net3 IN3 net1 VDD p12 l = 0.1u w = 0.35u m = 1
mmp3 net3 IN4 net1 VDD p12 l = 0.1u w = 0.35u m = 1
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp6 QN net5 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmn5 net5 net3 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net4 IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net3 IN3 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 QN net5 VSS VSS n12 l = 0.1u w = 0.43u m = 1


.ends AOI22X1



.subckt AOI22X2 IN1 IN2 IN3 IN4 QN VDD VSS
mmp4 net3 IN3 net1 VDD p12 l = 0.1u w = 0.35u m = 1
mmp6 QN net5 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp5 net5 net3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp3 net3 IN4 net1 VDD p12 l = 0.1u w = 0.35u m = 1
mmp1 net1 IN2 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmn6 QN net5 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn2 net3 IN1 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 net3 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn3 net4 IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net3 IN3 net4 VSS n12 l = 0.1u w = 0.21u m = 1


.ends AOI22X2



.subckt AOINVX1 INP VDD VDDG VSS ZN
mmn1 ZN INP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp1 ZN INP VDDG VDDG p12 l = 0.1u w = 0.5u m = 1


.ends AOINVX1



.subckt AOINVX2 INP VDD VDDG VSS ZN
mmn1 ZN INP VSS VSS n12 l = 0.1u w = 0.25u m = 2
mmp1 ZN INP VDDG VDDG p12 l = 0.1u w = 0.56u m = 2


.ends AOINVX2



.subckt AOINVX4 INP VDD VDDG VSS ZN
mmp1 ZN INP VDDG VDDG p12 l = 0.1u w = 1.12u m = 4
mmn1 ZN INP VSS VSS n12 l = 0.1u w = 0.49u m = 4


.ends AOINVX4



.subckt BSLEX1 ENB INOUT1 INOUT2 VDD VSS
mmn1 net1 ENB VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn2 INOUT1 ENB INOUT2 VSS n12 l = 0.1u w = 0.31u m = 1
mmp1 net1 ENB VDD VDD p12 l = 0.1u w = 0.28u m = 1
mmp2 INOUT1 net1 INOUT2 VDD p12 l = 0.1u w = 1.12u m = 1


.ends BSLEX1



.subckt BSLEX2 ENB INOUT1 INOUT2 VDD VSS
mmp2 INOUT1 net1 INOUT2 VDD p12 l = 0.1u w = 1.12u m = 2
mmp1 net1 ENB VDD VDD p12 l = 0.1u w = 0.56u m = 1

mmn1 net1 ENB VSS VSS n12 l = 0.1u w = 0.28u m = 1
mmn2 INOUT1 ENB INOUT2 VSS n12 l = 0.1u w = 0.31u m = 2

.ends BSLEX2



.subckt BSLEX4 ENB INOUT1 INOUT2 VDD VSS
mmp2 INOUT1 net1 INOUT2 VDD p12 l = 0.1u w = 1.12u m = 4
mmp1 net1 ENB VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmn1 net1 ENB VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn2 INOUT1 ENB INOUT2 VSS n12 l = 0.1u w = 0.31u m = 4


.ends BSLEX4



.subckt BUSKP INP VDD VSS
mg_nmos4t1 n3 net1 VSS VSS n12 l = 0.35u w = 0.21u m = 1
mg_nmos4t2 INP net1 n3 VSS n12 l = 0.35u w = 0.21u m = 1
mg_nmos4t3 net1 INP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mg_pmos4t1 n2 net1 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mg_pmos4t2 INP net1 n2 VDD p12 l = 0.1u w = 0.21u m = 1
mP1 net1 INP VDD VDD p12 l = 0.1u w = 0.65u m = 1


.ends BUSKP



.subckt CGLNPRX2 CLK EN GCLK SE VDD VSS
mmp12 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net3 CLKP net4 VDD p12 l = 0.1u w = 0.21u m = 1
mmp7 net6 ENL VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp11 CLKN CLK VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp2 net2 EN net1 VDD p12 l = 0.1u w = 0.21u m = 1
mmp3 net2 CLKN net3 VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 GCLK net7 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp4 ENL net3 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp8 net8 CLKP VDD VDD p12 l = 0.1u w = 0.58u m = 1
mmp5 net4 ENL VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net7 net6 net8 VDD p12 l = 0.1u w = 0.58u m = 1
mmp1 net1 SE VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmn11 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net5 ENL VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 GCLK net7 VSS VSS n12 l = 0.1u w = 0.53u m = 2
mmn3 net2 CLKP net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net7 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net3 CLKN net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 EN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 ENL net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net6 ENL VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn9 net7 net6 VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends CGLNPRX2



.subckt CGLNPRX8 CLK EN GCLK SE VDD VSS
mmn03 net2 CLKP net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net2 EN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 ENL net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net3 CLKN net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn06 net5 ENL VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 net2 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 GCLK net7 VSS VSS n12 l = 0.1u w = 0.56u m = 8
mmn09 net7 net6 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn08 net7 CLKP VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn07 net6 ENL VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmp03 net2 CLKN net3 VDD p12 l = 0.1u w = 0.21u m = 1
mmp01 net1 SE VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp11 CLKN CLK VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp04 ENL net3 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp06 net3 CLKP net4 VDD p12 l = 0.1u w = 0.21u m = 1
mmp05 net4 ENL VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp02 net2 EN net1 VDD p12 l = 0.1u w = 0.21u m = 1
mmp08 net8 CLKP VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp10 GCLK net7 VDD VDD p12 l = 0.1u w = 1.12u m = 8
mmp09 net7 net6 net8 VDD p12 l = 0.1u w = 1.12u m = 1
mmp07 net6 ENL VDD VDD p12 l = 0.1u w = 0.21u m = 1


.ends CGLNPRX8



.subckt CGLNPSX16 CLK EN GCLK SE VDD VSS
mmn4 net2 CLKN net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 ENL SE VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn12 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 CLKP VSS VSS n12 l = 0.1u w = 0.4u m = 2
mmn5 net4 net5 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net5 net2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 EN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net1 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net9 ENL VSS VSS n12 l = 0.1u w = 0.4u m = 2
mmn7 ENL net5 VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn11 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 GCLK net9 VSS VSS n12 l = 0.1u w = 0.475u m = 16
mmp4 net3 net5 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 net2 CLKP net3 VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 GCLK net9 VDD VDD p12 l = 0.1u w = 1.12u m = 16
mmp12 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp8 net8 CLKP VDD VDD p12 l = 0.1u w = 1.17u m = 2
mmp11 CLKN CLK VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp7 ENL net5 net6 VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net1 CLKN net2 VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net6 SE VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 EN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp3 net5 net2 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net9 ENL net8 VDD p12 l = 0.1u w = 1.17u m = 2


.ends CGLNPSX16



.subckt CGLNPSX2 CLK EN GCLK SE VDD VSS
mmn4 net2 CLKN net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 GCLK net9 VSS VSS n12 l = 0.1u w = 0.42u m = 2
mmn5 net4 net5 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net5 net2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 ENL SE VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn7 ENL net5 VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn1 net1 EN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net9 ENL VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net1 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmp7 ENL net5 net6 VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 GCLK net9 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp11 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 EN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net9 ENL net8 VDD p12 l = 0.1u w = 0.86u m = 1
mmp12 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net3 net5 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net1 CLKN net2 VDD p12 l = 0.1u w = 0.21u m = 1
mmp8 net8 CLKP VDD VDD p12 l = 0.1u w = 0.86u m = 1
mmp5 net2 CLKP net3 VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net6 SE VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp3 net5 net2 VDD VDD p12 l = 0.1u w = 0.21u m = 1


.ends CGLNPSX2



.subckt CGLNPSX4 CLK EN GCLK SE VDD VSS
mmn10 GCLK net9 VSS VSS n12 l = 0.1u w = 0.5u m = 4
mmn3 net5 net2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net1 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net2 CLKN net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 EN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net4 net5 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 ENL SE VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn9 net9 ENL VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 ENL net5 VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn8 net9 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp7 ENL net5 net6 VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 net2 CLKP net3 VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp11 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net6 SE VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 EN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp8 net8 CLKP VDD VDD p12 l = 0.1u w = 0.88u m = 1
mmp4 net3 net5 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net1 CLKN net2 VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 GCLK net9 VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmp3 net5 net2 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net9 ENL net8 VDD p12 l = 0.1u w = 0.88u m = 1


.ends CGLNPSX4



.subckt CGLNPSX8 CLK EN GCLK SE VDD VSS
mmn10 GCLK net9 VSS VSS n12 l = 0.1u w = 0.56u m = 8
mmn3 net5 net2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net1 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net2 CLKN net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 EN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net4 net5 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 ENL SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net9 ENL VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 ENL net5 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp7 ENL net5 net6 VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 net2 CLKP net3 VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp11 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net6 SE VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 EN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp8 net8 CLKP VDD VDD p12 l = 0.1u w = 0.9u m = 1
mmp4 net3 net5 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net1 CLKN net2 VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 GCLK net9 VDD VDD p12 l = 0.1u w = 1.12u m = 8
mmp3 net5 net2 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net9 ENL net8 VDD p12 l = 0.1u w = 0.9u m = 1


.ends CGLNPSX8



.subckt CGLPPRX2 CLK EN GCLK SE VDD VSS
mmn03 net2 CLKN net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net2 EN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 ENL net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net3 CLKP net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn06 net5 ENL VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 net2 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn07 net6 ENL net7 VSS n12 l = 0.1u w = 0.21u m = 1
mmn08 net7 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn09 GCLK net6 VSS VSS n12 l = 0.1u w = 0.53u m = 2
mmp03 net2 CLKP net3 VDD p12 l = 0.1u w = 0.21u m = 1
mmp01 net1 SE VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp11 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 CLKN CLK VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp04 ENL net3 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp06 net3 CLKN net4 VDD p12 l = 0.1u w = 0.21u m = 1
mmp05 net4 ENL VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp02 net2 EN net1 VDD p12 l = 0.1u w = 0.21u m = 1
mmp07 net6 ENL VDD VDD p12 l = 0.1u w = 0.24u m = 1
mmp08 net6 CLKP VDD VDD p12 l = 0.1u w = 0.24u m = 1
mmp09 GCLK net6 VDD VDD p12 l = 0.1u w = 1.12u m = 2


.ends CGLPPRX2



.subckt CGLPPRX8 CLK EN GCLK SE VDD VSS
mmn6 net5 ENL VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 EN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net6 ENL net7 VSS n12 l = 0.1u w = 0.68u m = 1
mmn1 net2 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 GCLK net6 VSS VSS n12 l = 0.1u w = 0.5u m = 8
mmn11 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn8 net7 CLKP VSS VSS n12 l = 0.1u w = 0.68u m = 1
mmn5 net3 CLKP net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 ENL net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 CLKN net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp11 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 ENL net3 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 net4 ENL VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 GCLK net6 VDD VDD p12 l = 0.1u w = 1.12u m = 8
mmp10 CLKN CLK VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp7 net6 ENL VDD VDD p12 l = 0.1u w = 0.87u m = 1
mmp8 net6 CLKP VDD VDD p12 l = 0.1u w = 0.87u m = 1
mmp2 net2 EN net1 VDD p12 l = 0.1u w = 0.21u m = 1
mmp3 net2 CLKP net3 VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 SE VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net3 CLKN net4 VDD p12 l = 0.1u w = 0.21u m = 1


.ends CGLPPRX8



.subckt CGLPPSX16 CLK EN GCLK SE VDD VSS
mmn9 net8 ENL net9 VSS n12 l = 0.1u w = 1.38u m = 1
mmn11 GCLK net8 VSS VSS n12 l = 0.1u w = 0.56u m = 16
mmn1 net1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 EN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net4 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 ENL net1 net7 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net3 CLKP net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net6 net4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net7 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net9 CLKP VSS VSS n12 l = 0.1u w = 1.38u m = 1
mmn13 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 CLKN net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp6 net3 CLKN net5 VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net2 EN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp8 ENL net3 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 net5 net4 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 SE VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp7 ENL net1 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net8 CLKP VDD VDD p12 l = 0.1u w = 0.32u m = 4
mmp12 CLKN CLK VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp4 net4 net3 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp3 net2 CLKP net3 VDD p12 l = 0.1u w = 0.21u m = 1
mmp11 GCLK net8 VDD VDD p12 l = 0.1u w = 1.12u m = 16
mmp9 net8 ENL VDD VDD p12 l = 0.1u w = 0.32u m = 4


.ends CGLPPSX16



.subckt CGLPPSX2 CLK EN GCLK SE VDD VSS
mmn03 net2 CLKN net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn07 ENL net1 net7 VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 net4 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net3 CLKP net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn06 net6 net4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn08 net7 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn09 net8 ENL net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net9 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 GCLK net8 VSS VSS n12 l = 0.1u w = 0.56u m = 2
mmn01 net1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net2 EN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp03 net2 CLKP net3 VDD p12 l = 0.1u w = 0.21u m = 1
mmp07 ENL net1 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 CLKN CLK VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp04 net4 net3 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp06 net3 CLKN net5 VDD p12 l = 0.1u w = 0.21u m = 1
mmp05 net5 net4 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp08 ENL net3 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp09 net8 ENL VDD VDD p12 l = 0.1u w = 0.24u m = 1
mmp10 net8 CLKP VDD VDD p12 l = 0.1u w = 0.24u m = 1
mmp11 GCLK net8 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp01 net1 SE VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp02 net2 EN VDD VDD p12 l = 0.1u w = 0.21u m = 1


.ends CGLPPSX2



.subckt CGLPPSX4 CLK EN GCLK SE VDD VSS
mmp13 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 ENL VDD VDD p12 l = 0.1u w = 0.28u m = 1
mmp7 ENL net1 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net3 CLKN net5 VDD p12 l = 0.1u w = 0.21u m = 1
mmp3 net2 CLKP net3 VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net8 CLKP VDD VDD p12 l = 0.1u w = 0.28u m = 1
mmp11 GCLK net8 VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmp2 net2 EN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 net5 net4 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net4 net3 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp8 ENL net3 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 SE VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 CLKN CLK VDD VDD p12 l = 0.1u w = 0.42u m = 1

mmn12 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 ENL net1 net7 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 EN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net4 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 ENL net9 VSS n12 l = 0.1u w = 0.25u m = 1
mmn1 net1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 CLKN net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net6 net4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 GCLK net8 VSS VSS n12 l = 0.1u w = 0.56u m = 4
mmn13 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.41u m = 1
mmn8 net7 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net9 CLKP VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn5 net3 CLKP net6 VSS n12 l = 0.1u w = 0.21u m = 1

.ends CGLPPSX4



.subckt CGLPPSX8 CLK EN GCLK SE VDD VSS
mmn13 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 GCLK net8 VSS VSS n12 l = 0.1u w = 0.55u m = 8
mmn6 net6 net4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 CLKN net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net9 CLKP VSS VSS n12 l = 0.1u w = 0.69u m = 1
mmn9 net8 ENL net9 VSS n12 l = 0.1u w = 0.69u m = 1
mmn8 net7 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net3 CLKP net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 EN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 ENL net1 net7 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net4 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp12 CLKN CLK VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp2 net2 EN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp11 GCLK net8 VDD VDD p12 l = 0.1u w = 1.12u m = 8
mmp9 net8 ENL VDD VDD p12 l = 0.1u w = 0.7u m = 1
mmp1 net1 SE VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net3 CLKN net5 VDD p12 l = 0.1u w = 0.21u m = 1
mmp3 net2 CLKP net3 VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 net5 net4 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp8 ENL net3 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net4 net3 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp7 ENL net1 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net8 CLKP VDD VDD p12 l = 0.1u w = 0.7u m = 1
mmp13 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1


.ends CGLPPSX8



.subckt CLOAD1 INP VDD VSS
mmp1 VDD INP VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmn1 VSS INP VSS VSS n12 l = 0.1u w = 0.49u m = 1


.ends CLOAD1



.subckt DCAP VDD VSS
mg_nmos4t1 _n1 _n6 VSS VSS n12 l = 0.1u w = 0.69u m = 1
mg_pmos4t1 _n6 _n1 VDD VDD p12 l = 0.1u w = 0.8u m = 1


.ends DCAP



.subckt DEC24X1 IN1 IN2 Q0 Q1 Q2 Q3 VDD VSS
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.41u m = 1
mmp3 net3 net1 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp6 net4 IN2 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp2 net2 IN2 VDD VDD p12 l = 0.1u w = 0.41u m = 1
mmp5 net4 net1 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp12 Q1 net4 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp7 net5 IN1 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp8 net5 net2 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp9 net6 IN1 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp10 net6 IN2 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp11 Q0 net3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp4 net3 net2 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp13 Q2 net5 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp14 Q3 net6 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmn1 net1 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 _n10 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 Q0 net3 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net4 IN2 _n130 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 _n130 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net5 net2 _n148 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 _n148 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net6 IN2 _n166 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 _n166 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net3 net2 _n10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 Q1 net4 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn13 Q2 net5 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn14 Q3 net6 VSS VSS n12 l = 0.1u w = 0.4u m = 1


.ends DEC24X1



.subckt DEC24X2 IN1 IN2 Q0 Q1 Q2 Q3 VDD VSS
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp3 net3 net1 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp6 net4 IN2 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp2 net2 IN2 VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp5 net4 net1 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp12 Q1 net4 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp7 net5 IN1 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp8 net5 net2 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp9 net6 IN1 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp10 net6 IN2 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp11 Q0 net3 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp4 net3 net2 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp13 Q2 net5 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp14 Q3 net6 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmn1 net1 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 _n10 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 Q0 net3 VSS VSS n12 l = 0.1u w = 0.4u m = 2
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net4 IN2 _n130 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 _n130 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net5 net2 _n148 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 _n148 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net6 IN2 _n166 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 _n166 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net3 net2 _n10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 Q1 net4 VSS VSS n12 l = 0.1u w = 0.4u m = 2
mmn13 Q2 net5 VSS VSS n12 l = 0.1u w = 0.4u m = 2
mmn14 Q3 net6 VSS VSS n12 l = 0.1u w = 0.4u m = 2


.ends DEC24X2



.subckt DELLN1X2 INP VDD VSS Z
mmp1 net1 INP VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net01 VSS VDD VDD p12 l = 0.1u w = 0.2u m = 1
mmp3 net2 net1 net01 VDD p12 l = 0.1u w = 0.2u m = 1
mmp4 net3 net2 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 Z net3 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmn3 net2 net1 net02 VSS n12 l = 0.2u w = 0.14u m = 1
mmn2 net02 VDD VSS VSS n12 l = 0.2u w = 0.14u m = 1
mmn1 net1 INP VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn5 Z net3 VSS VSS n12 l = 0.1u w = 0.41u m = 2
mmn4 net3 net2 VSS VSS n12 l = 0.2u w = 0.14u m = 1


.ends DELLN1X2



.subckt DELLN2X2 INP VDD VSS Z
mmp1 net1 INP VDD VDD p12 l = 0.1u w = 0.14u m = 1
mmp2 net01 VSS VDD VDD p12 l = 0.13u w = 0.14u m = 1
mmp3 net2 net1 net01 VDD p12 l = 0.13u w = 0.14u m = 1
mmp4 net3 net2 VDD VDD p12 l = 0.14u w = 0.15u m = 1
mmp5 Z net3 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmn3 net2 net1 net02 VSS n12 l = 0.37u w = 0.14u m = 1
mmn2 net02 VDD VSS VSS n12 l = 0.37u w = 0.14u m = 1
mmn1 net1 INP VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn5 Z net3 VSS VSS n12 l = 0.1u w = 0.42u m = 2
mmn4 net3 net2 VSS VSS n12 l = 0.37u w = 0.14u m = 1


.ends DELLN2X2



.subckt DELLN3X2 INP VDD VSS Z
mmp1 net1 INP VDD VDD p12 l = 0.1u w = 0.14u m = 1
mmp2 net01 VSS VDD VDD p12 l = 0.12u w = 0.14u m = 1
mmp3 net2 net1 net01 VDD p12 l = 0.12u w = 0.14u m = 1
mmp6 net4 net3 net03 VDD p12 l = 0.12u w = 0.14u m = 1
mmp5 net03 VSS VDD VDD p12 l = 0.12u w = 0.14u m = 1
mmp7 net5 net4 VDD VDD p12 l = 0.11u w = 0.14u m = 1
mmp4 net3 net2 VDD VDD p12 l = 0.12u w = 0.14u m = 1
mmp8 Z net5 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmn6 net4 net3 net04 VSS n12 l = 0.36u w = 0.14u m = 1
mmn5 net04 VDD VSS VSS n12 l = 0.36u w = 0.14u m = 1
mmn3 net2 net1 net02 VSS n12 l = 0.36u w = 0.14u m = 1
mmn2 net02 VDD VSS VSS n12 l = 0.36u w = 0.14u m = 1
mmn1 net1 INP VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn7 net5 net4 VSS VSS n12 l = 0.29u w = 0.14u m = 1
mmn8 Z net5 VSS VSS n12 l = 0.1u w = 0.42u m = 2
mmn4 net3 net2 VSS VSS n12 l = 0.36u w = 0.14u m = 1


.ends DELLN3X2



.subckt DFFARX1 CLK D Q QN RSTB VDD VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.44u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.52u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFARX1



.subckt DFFARX2 CLK D Q QN RSTB VDD VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.2u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.76u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFARX2



.subckt DFFASRX1 CLK D Q QN RSTB SETB VDD VSS
mmp01 net01 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.3u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKP net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 net01 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net01 VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFASRX1



.subckt DFFASRX2 CLK D Q QN RSTB SETB VDD VSS
mmp01 net01 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKP net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 net01 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 1.1u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.8u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net01 VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFASRX2



.subckt DFFASX1 CLK D Q QN SETB VDD VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.45u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFASX1



.subckt DFFASX2 CLK D Q QN SETB VDD VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.53u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.2u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFASX2



.subckt DFFNARX1 CLK D Q QN RSTB VDD VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 0.9u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.5u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.32u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.32u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.35u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFNARX1



.subckt DFFNARX2 CLK D Q QN RSTB VDD VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp1 net1 CLKN net06 VDD p12 l = 0.1u w = 0.5u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.5u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.6u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFNARX2



.subckt DFFNASRNX1 CLK D QN RSTB SETB VDD VSS
mmp01 net01 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKN net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 net01 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.53u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net01 VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFNASRNX1



.subckt DFFNASRNX2 CLK D QN RSTB SETB VDD VSS
mmp01 net01 D VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.5u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKN net01 VDD p12 l = 0.1u w = 0.5u m = 1
mmn01 net01 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 1.1u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net01 VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFNASRNX2



.subckt DFFNASRQX1 CLK D Q RSTB SETB VDD VSS
mmp01 net01 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.26u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKN net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 net01 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.48u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net01 VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFNASRQX1



.subckt DFFNASRQX2 CLK D Q RSTB SETB VDD VSS
mmp01 net01 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKN net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 net01 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.7u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net01 VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFNASRQX2



.subckt DFFNASRX1 CLK D Q QN RSTB SETB VDD VSS
mmp01 net01 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKN net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 net01 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.48u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.48u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net01 VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFNASRX1



.subckt DFFNASRX2 CLK D Q QN RSTB SETB VDD VSS
mmp01 net22 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKN net22 VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 net22 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 1.1u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.7u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net22 VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFNASRX2



.subckt DFFNASX1 CLK D Q QN SETB VDD VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.37u m = 1
mmp1 net1 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.45u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.52u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFNASX1



.subckt DFFNASX2 CLK D Q QN SETB VDD VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.53u m = 1
mmp1 net1 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.2u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFNASX2



.subckt DFFNX1 CLK D Q QN VDD VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.5u m = 1
mmp1 net1 CLKN net06 VDD p12 l = 0.1u w = 0.5u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.4u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFNX1



.subckt DFFNX2 CLK D Q QN VDD VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.6u m = 1
mmp1 net1 CLKN net06 VDD p12 l = 0.1u w = 0.6u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.4u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.6u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFNX2



.subckt DFFSSRX1 CLK D Q QN RSTB SETB VDD VSS
mmp03 net06 D net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 net01 SET VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net06 RSTB net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN IQN VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp12 IQN net8 net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp8 net8 IQN VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 IQN CLKN net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp01 SET SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 net03 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 SET net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN IQN VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 IQN net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 IQN VSS VSS n12 l = 0.1u w = 0.35u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 IQN CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn01 SET SETB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFSSRX1



.subckt DFFSSRX2 CLK D Q QN RSTB SETB VDD VSS
mmp03 net06 D net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 net01 SET VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net06 RSTB net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN IQN VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp12 IQN net8 net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp8 net8 IQN VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 IQN CLKN net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp01 SET SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 net03 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 SET net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN IQN VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 IQN net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 IQN VSS VSS n12 l = 0.1u w = 0.35u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 IQN CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 1u m = 1
mmn01 SET SETB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFSSRX2



.subckt DFFX1 CLK D Q QN VDD VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFX1



.subckt DFFX2 CLK D Q QN VDD VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.56u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends DFFX2



.subckt DHFILLHLH2 VDD VSS


.ends DHFILLHLH2



.subckt DHFILLHLHLS11 VDDH VDDL VSS


.ends DHFILLHLHLS11



.subckt DHFILLLHL2 VDD VSS


.ends DHFILLLHL2



.subckt FADDX1 A B CI CO S VDD VSS
mmp2 net1 B VDD VDD p12 l = 0.1u w = 0.89u m = 1
mmp1 net1 A VDD VDD p12 l = 0.1u w = 0.89u m = 1
mmp5 net3 B net4 VDD p12 l = 0.1u w = 0.89u m = 1
mmp4 net4 A VDD VDD p12 l = 0.1u w = 0.89u m = 1
mmp7 net6 A VDD VDD p12 l = 0.1u w = 0.89u m = 1
mmp6 net6 CI VDD VDD p12 l = 0.1u w = 0.89u m = 1
mmp3 net3 CI net1 VDD p12 l = 0.1u w = 0.89u m = 1
mmp8 net6 B VDD VDD p12 l = 0.1u w = 0.89u m = 1
mmp9 net8 net3 net6 VDD p12 l = 0.1u w = 0.89u m = 1
mmp10 net9 A VDD VDD p12 l = 0.1u w = 0.89u m = 1
mmp11 net10 B net9 VDD p12 l = 0.1u w = 0.89u m = 1
mmp12 net8 CI net10 VDD p12 l = 0.1u w = 0.89u m = 1
mmp13 S net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp14 CO net3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmn5 net5 A VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn7 net7 A VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn4 net3 B net5 VSS n12 l = 0.1u w = 0.3u m = 1
mmn6 net7 CI VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn3 net2 B VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn2 net3 CI net2 VSS n12 l = 0.1u w = 0.3u m = 1
mmn1 net2 A VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn8 net8 net3 net7 VSS n12 l = 0.1u w = 0.3u m = 1
mmn9 net7 B VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn10 net8 CI net11 VSS n12 l = 0.1u w = 0.3u m = 1
mmn11 net11 B net12 VSS n12 l = 0.1u w = 0.3u m = 1
mmn12 net12 A VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn13 S net8 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn14 CO net3 VSS VSS n12 l = 0.1u w = 0.48u m = 1


.ends FADDX1



.subckt FADDX2 A B CI CO S VDD VSS
mmp2 net1 B VDD VDD p12 l = 0.1u w = 0.89u m = 1
mmp1 net1 A VDD VDD p12 l = 0.1u w = 0.89u m = 1
mmp5 net3 B net4 VDD p12 l = 0.1u w = 0.89u m = 1
mmp4 net4 A VDD VDD p12 l = 0.1u w = 0.89u m = 1
mmp7 net6 A VDD VDD p12 l = 0.1u w = 0.89u m = 1
mmp6 net6 CI VDD VDD p12 l = 0.1u w = 0.89u m = 1
mmp3 net3 CI net1 VDD p12 l = 0.1u w = 0.89u m = 1
mmp8 net6 B VDD VDD p12 l = 0.1u w = 0.89u m = 1
mmp9 net8 net3 net6 VDD p12 l = 0.1u w = 0.89u m = 1
mmp10 net9 A VDD VDD p12 l = 0.1u w = 0.89u m = 1
mmp11 net10 B net9 VDD p12 l = 0.1u w = 0.89u m = 1
mmp12 net8 CI net10 VDD p12 l = 0.1u w = 0.89u m = 1
mmp13 S net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp14 CO net3 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmn5 net5 A VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn7 net7 A VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn4 net3 B net5 VSS n12 l = 0.1u w = 0.3u m = 1
mmn6 net7 CI VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn3 net2 B VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn2 net3 CI net2 VSS n12 l = 0.1u w = 0.3u m = 1
mmn1 net2 A VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn8 net8 net3 net7 VSS n12 l = 0.1u w = 0.3u m = 1
mmn9 net7 B VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn10 net8 CI net11 VSS n12 l = 0.1u w = 0.3u m = 1
mmn11 net11 B net12 VSS n12 l = 0.1u w = 0.3u m = 1
mmn12 net12 A VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn13 S net8 VSS VSS n12 l = 0.1u w = 1u m = 1
mmn14 CO net3 VSS VSS n12 l = 0.1u w = 0.96u m = 1


.ends FADDX2



.subckt HADDX1 A0 B0 C1 SO VDD VSS
mmp3 net2 net4 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp2 net2 B0 net1 VDD p12 l = 0.1u w = 0.7u m = 1
mmp1 net1 A0 VDD VDD p12 l = 0.1u w = 0.7u m = 1
mmp4 net4 A0 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp5 net4 B0 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp6 SO net2 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp7 C1 net4 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmn1 net2 A0 net3 VSS n12 l = 0.1u w = 0.3u m = 1
mmn3 net3 net4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 SO net2 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn4 net5 A0 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net4 B0 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 B0 net3 VSS n12 l = 0.1u w = 0.3u m = 1
mmn7 C1 net4 VSS VSS n12 l = 0.1u w = 0.4u m = 1


.ends HADDX1



.subckt HADDX2 A0 B0 C1 SO VDD VSS
mmp3 net2 net4 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp2 net2 B0 net1 VDD p12 l = 0.1u w = 0.7u m = 1
mmp1 net1 A0 VDD VDD p12 l = 0.1u w = 0.7u m = 1
mmp4 net4 A0 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp5 net4 B0 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp6 SO net2 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp7 C1 net4 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmn1 net2 A0 net3 VSS n12 l = 0.1u w = 0.3u m = 1
mmn3 net3 net4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 SO net2 VSS VSS n12 l = 0.1u w = 0.4u m = 2
mmn4 net5 A0 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net4 B0 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 B0 net3 VSS n12 l = 0.1u w = 0.3u m = 1
mmn7 C1 net4 VSS VSS n12 l = 0.1u w = 0.4u m = 2


.ends HADDX2



.subckt HEAD2X16 SLEEP SLEEPOUT VDD VDDG VSS


mg_pmos4t_hvt1 VDD net0 VDDG VDDG p12_hvt l = 0.1u w = 1.12u m = 16
mg_nmos4t2 SLEEPOUT net0 VDDG VDDG p12 l = 0.1u w = 1.1u m = 16
mg_nmos4t1 net0 SLEEP VDDG VDDG p12 l = 0.1u w = 0.48u m = 1
mg_pmos4t2 SLEEPOUT net0 VSS VSS n12 l = 0.1u w = 0.49u m = 16
mg_pmos4t1 net0 SLEEP VSS VSS n12 l = 0.1u w = 0.24u m = 1
.ends HEAD2X16



.subckt HEAD2X2 SLEEP SLEEPOUT VDD VDDG VSS

mg_pmos4t_hvt1 VDD net0 VDDG VDDG p12_hvt l = 0.1u w = 2.24u m = 1
mg_pmos4t1 net0 SLEEP VSS VSS n12 l = 0.1u w = 0.24u m = 1
mg_pmos4t2 SLEEPOUT net0 VSS VSS n12 l = 0.1u w = 0.49u m = 2
mg_nmos4t2 SLEEPOUT net0 VDDG VDDG p12 l = 0.1u w = 1.12u m = 2
mg_nmos4t1 net0 SLEEP VDDG VDDG p12 l = 0.1u w = 0.48u m = 1

.ends HEAD2X2



.subckt HEAD2X32 SLEEP SLEEPOUT VDD VDDG VSS


mg_pmos4t_hvt1 VDD net0 VDDG VDDG p12_hvt l = 0.1u w = 1.12u m = 32
mg_nmos4t2 SLEEPOUT net0 VDDG VDDG p12 l = 0.1u w = 1.1u m = 32
mg_nmos4t1 net0 SLEEP VDDG VDDG p12 l = 0.1u w = 0.48u m = 1
mg_pmos4t2 SLEEPOUT net0 VSS VSS n12 l = 0.1u w = 0.49u m = 32
mg_pmos4t1 net0 SLEEP VSS VSS n12 l = 0.1u w = 0.24u m = 1
.ends HEAD2X32



.subckt HEAD2X4 SLEEP SLEEPOUT VDD VDDG VSS
mg_pmos4t3 VDD net0 VDDG VDDG p12_hvt l = 0.1u w = 1.12u m = 4


mg_pmos4t1 net0 SLEEP VDDG VDDG p12 l = 0.1u w = 0.5u m = 1
mg_pmos4t2 SLEEPOUT net0 VDDG VDDG p12 l = 0.1u w = 1.1u m = 4
mg_nmos4t2 SLEEPOUT net0 VSS VSS n12 l = 0.1u w = 0.49u m = 4
mg_nmos4t1 net0 SLEEP VSS VSS n12 l = 0.1u w = 0.24u m = 1
.ends HEAD2X4



.subckt HEAD2X8 SLEEP SLEEPOUT VDD VDDG VSS


mg_pmos4t_hvt1 VDD net0 VDDG VDDG p12_hvt l = 0.1u w = 1.12u m = 8
mg_nmos4t2 SLEEPOUT net0 VDDG VDDG p12 l = 0.1u w = 1.1u m = 8
mg_nmos4t1 net0 SLEEP VDDG VDDG p12 l = 0.1u w = 0.48u m = 1
mg_pmos4t2 SLEEPOUT net0 VSS VSS n12 l = 0.1u w = 0.49u m = 8
mg_pmos4t1 net0 SLEEP VSS VSS n12 l = 0.1u w = 0.24u m = 1
.ends HEAD2X8



.subckt HEADX16 SLEEP VDD VDDG VSS


mg_pmos4t_hvt1 VDD SLEEP VDDG VDDG p12_hvt l = 0.1u w = 1.12u m = 16
.ends HEADX16



.subckt HEADX2 SLEEP VDD VDDG VSS


mg_pmos4t_hvt1 VDD SLEEP VDDG VDDG p12_hvt l = 0.1u w = 2.24u m = 1
.ends HEADX2



.subckt HEADX32 SLEEP VDD VDDG VSS


mg_pmos4t_hvt1 VDD SLEEP VDDG VDDG p12_hvt l = 0.1u w = 1.12u m = 32
.ends HEADX32



.subckt HEADX4 SLEEP VDD VDDG VSS


mg_pmos4t_hvt1 VDD SLEEP VDDG VDDG p12_hvt l = 0.1u w = 1.12u m = 4
.ends HEADX4



.subckt HEADX8 SLEEP VDD VDDG VSS


mg_pmos4t_hvt1 VDD SLEEP VDDG VDDG p12_hvt l = 0.1u w = 1.12u m = 8
.ends HEADX8



.subckt IBUFFX16 INP VDD VSS ZN

mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp3 ZN net2 VDD VDD p12 l = 0.1u w = 1.12u m = 16
mmp1 net1 INP VDD VDD p12 l = 0.1u w = 0.5u m = 1

mmn3 ZN net2 VSS VSS n12 l = 0.1u w = 0.43u m = 16
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn1 net1 INP VSS VSS n12 l = 0.1u w = 0.21u m = 1
.ends IBUFFX16



.subckt IBUFFX2 INP VDD VSS ZN
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.62u m = 1
mmp3 ZN net2 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp1 net1 INP VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmn3 ZN net2 VSS VSS n12 l = 0.1u w = 0.45u m = 2
mmn1 net1 INP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends IBUFFX2



.subckt IBUFFX32 INP VDD VSS ZN
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmp3 ZN net2 VDD VDD p12 l = 0.1u w = 1.12u m = 32
mmp1 net1 INP VDD VDD p12 l = 0.1u w = 0.5u m = 1

mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.43u m = 4
mmn3 ZN net2 VSS VSS n12 l = 0.1u w = 0.43u m = 32
mmn1 net1 INP VSS VSS n12 l = 0.1u w = 0.21u m = 1

.ends IBUFFX32



.subckt IBUFFX4 INP VDD VSS ZN
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp3 ZN net2 VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmp1 net1 INP VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmn3 ZN net2 VSS VSS n12 l = 0.1u w = 0.43u m = 4
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net1 INP VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends IBUFFX4



.subckt IBUFFX8 INP VDD VSS ZN
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp3 ZN net2 VDD VDD p12 l = 0.1u w = 1.12u m = 8
mmp1 net1 INP VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmn3 ZN net2 VSS VSS n12 l = 0.1u w = 0.43u m = 8
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net1 INP VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends IBUFFX8



.subckt INVX0 INP VDD VSS ZN
mmp1 ZN INP VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmn1 ZN INP VSS VSS n12 l = 0.1u w = 0.24u m = 1


.ends INVX0



.subckt INVX16 INP VDD VSS ZN
mmn1 ZN INP VSS VSS n12 l = 0.1u w = 0.49u m = 16
mmp1 ZN INP VDD VDD p12 l = 0.1u w = 1.12u m = 16


.ends INVX16



.subckt INVX1 INP VDD VSS ZN
mmp1 ZN INP VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmn1 ZN INP VSS VSS n12 l = 0.1u w = 0.49u m = 1


.ends INVX1



.subckt INVX2 INP VDD VSS ZN
mmp1 ZN INP VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmn1 ZN INP VSS VSS n12 l = 0.1u w = 0.49u m = 2


.ends INVX2



.subckt INVX32 INP VDD VSS ZN
mmn1 ZN INP VSS VSS n12 l = 0.1u w = 0.49u m = 32
mmp1 ZN INP VDD VDD p12 l = 0.1u w = 1.12u m = 32


.ends INVX32



.subckt INVX4 INP VDD VSS ZN
mmp1 ZN INP VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmn1 ZN INP VSS VSS n12 l = 0.1u w = 0.49u m = 4


.ends INVX4



.subckt INVX8 INP VDD VSS ZN
mmn1 ZN INP VSS VSS n12 l = 0.1u w = 0.49u m = 8
mmp1 ZN INP VDD VDD p12 l = 0.1u w = 1.12u m = 8


.ends INVX8



.subckt ISOLANDAOX1 D ISO Q VDD VDDG VSS
mmp3 outnand D VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp2 outnand ISON VDDG VDDG p12 l = 0.1u w = 0.31u m = 1
mmp4 Q outnand VDDG VDDG p12 l = 0.1u w = 1.1u m = 1
mmp1 ISON ISO VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmn3 outnand D netn2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 Q outnand VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn2 netn2 ISON VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 ISON ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends ISOLANDAOX1



.subckt ISOLANDAOX2 D ISO Q VDD VDDG VSS
mmp3 outnand D VDD VDD p12 l = 0.1u w = 0.37u m = 1
mmp2 outnand ISON VDDG VDDG p12 l = 0.1u w = 0.31u m = 1
mmp4 Q outnand VDDG VDDG p12 l = 0.1u w = 1.1u m = 2
mmp1 ISON ISO VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmn3 outnand D netn2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 Q outnand VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn2 netn2 ISON VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 ISON ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends ISOLANDAOX2



.subckt ISOLANDAOX4 D ISO Q VDD VDDG VSS
mmp3 outnand D VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp2 outnand ISON VDDG VDDG p12 l = 0.1u w = 0.31u m = 1
mmp4 Q outnand VDDG VDDG p12 l = 0.1u w = 1.1u m = 4
mmp1 ISON ISO VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmn3 outnand D netn2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 Q outnand VSS VSS n12 l = 0.1u w = 0.5u m = 4
mmn2 netn2 ISON VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 ISON ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends ISOLANDAOX4



.subckt ISOLANDAOX8 D ISO Q VDD VDDG VSS
mmp3 outnand D VDD VDD p12 l = 0.1u w = 0.7u m = 1
mmp2 outnand ISON VDDG VDDG p12 l = 0.1u w = 0.7u m = 1
mmp4 Q outnand VDDG VDDG p12 l = 0.1u w = 1.1u m = 8
mmp1 ISON ISO VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmn3 outnand D netn2 VSS n12 l = 0.1u w = 0.4u m = 1
mmn4 Q outnand VSS VSS n12 l = 0.1u w = 0.5u m = 8
mmn2 netn2 ISON VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn1 ISON ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends ISOLANDAOX8



.subckt ISOLANDX1 D ISO Q VDD VSS
mmp3 outnand D VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp2 outnand ISON VDD VDD p12 l = 0.1u w = 0.31u m = 1
mmp4 Q outnand VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp1 ISON ISO VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn3 outnand D netn2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 Q outnand VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn2 netn2 ISON VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 ISON ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends ISOLANDX1



.subckt ISOLANDX2 D ISO Q VDD VSS
mmp3 outnand D VDD VDD p12 l = 0.1u w = 0.37u m = 1
mmp2 outnand ISON VDD VDD p12 l = 0.1u w = 0.31u m = 1
mmp4 Q outnand VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp1 ISON ISO VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn3 outnand D netn2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 Q outnand VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn2 netn2 ISON VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 ISON ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends ISOLANDX2



.subckt ISOLANDX4 D ISO Q VDD VSS
mmp3 outnand D VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp2 outnand ISON VDD VDD p12 l = 0.1u w = 0.31u m = 1
mmp4 Q outnand VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmp1 ISON ISO VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn3 outnand D netn2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 Q outnand VSS VSS n12 l = 0.1u w = 0.5u m = 4
mmn2 netn2 ISON VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 ISON ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends ISOLANDX4



.subckt ISOLANDX8 D ISO Q VDD VSS
mmp3 outnand D VDD VDD p12 l = 0.1u w = 0.7u m = 1
mmp2 outnand ISON VDD VDD p12 l = 0.1u w = 0.7u m = 1
mmp4 Q outnand VDD VDD p12 l = 0.1u w = 1.12u m = 8
mmp1 ISON ISO VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn3 outnand D netn2 VSS n12 l = 0.1u w = 0.4u m = 1
mmn4 Q outnand VSS VSS n12 l = 0.1u w = 0.5u m = 8
mmn2 netn2 ISON VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn1 ISON ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends ISOLANDX8



.subckt ISOLORAOX1 D ISO Q VDD VDDG VSS
mmn1 netp2 ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 Q netp2 VSS VSS n12 l = 0.1u w = 0.48u m = 1
mmn2 netp2 a VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 a net1 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmp4 a net1 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp2 netp2 a netp1 VDDG p12 l = 0.1u w = 0.9u m = 1
mmp3 Q netp2 VDDG VDDG p12 l = 0.1u w = 1.12u m = 1
mmp1 netp1 ISO VDDG VDDG p12 l = 0.1u w = 0.9u m = 1
mmp5 net1 D VDD VDD p12 l = 0.1u w = 0.62u m = 1

.ends ISOLORAOX1



.subckt ISOLORAOX2 D ISO Q VDD VDDG VSS
mmn3 Q netp2 VSS VSS n12 l = 0.1u w = 0.48u m = 2
mmn2 netp2 a VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 a net1 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn4 net1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp4 a net1 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp2 netp2 a netp1 VDDG p12 l = 0.1u w = 0.9u m = 1
mmp3 Q netp2 VDDG VDDG p12 l = 0.1u w = 1.12u m = 2
mmp5 net1 D VDD VDD p12 l = 0.1u w = 0.62u m = 1
mmp1 netp1 ISO VDDG VDDG p12 l = 0.1u w = 0.9u m = 1

.ends ISOLORAOX2



.subckt ISOLORAOX4 D ISO Q VDD VDDG VSS
mmn4 netp2 a VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 Q netp2 VSS VSS n12 l = 0.1u w = 0.48u m = 4
mmn6 netp2 ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 a net1 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn8 net1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp4 Q netp2 VDDG VDDG p12 l = 0.1u w = 1.12u m = 4
mmp5 netp2 a netp1 VDDG p12 l = 0.1u w = 0.9u m = 1
mmp6 a net1 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp7 net1 D VDD VDD p12 l = 0.1u w = 0.62u m = 1
mmp8 netp1 ISO VDDG VDDG p12 l = 0.1u w = 0.9u m = 1

.ends ISOLORAOX4



.subckt ISOLORAOX8 D ISO Q VDD VDDG VSS
mmn5 Q netp2 VSS VSS n12 l = 0.1u w = 0.48u m = 8
mmn6 netp2 ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 a net1 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn8 net1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp2 a VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp7 net1 D VDD VDD p12 l = 0.1u w = 0.62u m = 1
mmp4 Q netp2 VDDG VDDG p12 l = 0.1u w = 1.12u m = 8
mmp8 netp1 ISO VDDG VDDG p12 l = 0.1u w = 0.9u m = 1
mmp5 netp2 a netp1 VDDG p12 l = 0.1u w = 0.9u m = 1
mmp6 a net1 VDD VDD p12 l = 0.1u w = 1.12u m = 2

.ends ISOLORAOX8



.subckt ISOLORX1 D ISO Q VDD VSS
mmn1 netp2 ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 Q netp2 VSS VSS n12 l = 0.1u w = 0.48u m = 1
mmn2 netp2 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 netp2 D netp1 VDD p12 l = 0.1u w = 0.9u m = 1
mmp3 Q netp2 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp1 netp1 ISO VDD VDD p12 l = 0.1u w = 0.9u m = 1


.ends ISOLORX1



.subckt ISOLORX2 D ISO Q VDD VSS
mmn1 netp2 ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 Q netp2 VSS VSS n12 l = 0.1u w = 0.48u m = 2
mmn2 netp2 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 netp2 D netp1 VDD p12 l = 0.1u w = 0.95u m = 1
mmp3 Q netp2 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp1 netp1 ISO VDD VDD p12 l = 0.1u w = 0.95u m = 1


.ends ISOLORX2



.subckt ISOLORX4 D ISO Q VDD VSS
mmn1 netp2 ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 Q netp2 VSS VSS n12 l = 0.1u w = 0.5u m = 4
mmn2 netp2 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 netp2 D netp1 VDD p12 l = 0.1u w = 0.9u m = 1
mmp3 Q netp2 VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmp1 netp1 ISO VDD VDD p12 l = 0.1u w = 0.9u m = 1


.ends ISOLORX4



.subckt ISOLORX8 D ISO Q VDD VSS
mmn1 netp2 ISO VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 Q netp2 VSS VSS n12 l = 0.1u w = 0.5u m = 8
mmn2 netp2 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 netp2 D netp1 VDD p12 l = 0.1u w = 1.12u m = 1
mmp3 Q netp2 VDD VDD p12 l = 0.1u w = 1.12u m = 8
mmp1 netp1 ISO VDD VDD p12 l = 0.1u w = 1.12u m = 1


.ends ISOLORX8



.subckt LARX1 CLK D Q QN RSTB VDD VSS
mmp5 net3 IQN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q net5 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp7 net5 net3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp9 QN net3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp2 net1 RSTB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 IQN CLKN net1 VDD p12 l = 0.1u w = 0.25u m = 1
mmp4 net5 CLKP IQN VDD p12 l = 0.1u w = 0.21u m = 1
mmp8 net5 RSTB VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmn1 net2 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net5 CLKN IQN VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q net5 VSS VSS n12 l = 0.1u w = 0.49u m = 1
mmn2 net1 RSTB net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net3 IQN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 QN net3 VSS VSS n12 l = 0.1u w = 0.49u m = 1
mmn8 net6 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net5 net3 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 IQN CLKP net1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends LARX1



.subckt LARX2 CLK D Q QN RSTB VDD VSS
mmp5 net3 IQN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q net5 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp7 net5 net3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp9 QN net3 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp2 net1 RSTB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 IQN CLKN net1 VDD p12 l = 0.1u w = 0.25u m = 1
mmp4 net5 CLKP IQN VDD p12 l = 0.1u w = 0.21u m = 1
mmp8 net5 RSTB VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmn1 net2 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net5 CLKN IQN VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q net5 VSS VSS n12 l = 0.1u w = 0.98u m = 1
mmn2 net1 RSTB net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net3 IQN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 QN net3 VSS VSS n12 l = 0.1u w = 0.98u m = 1
mmn8 net6 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net5 net3 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 IQN CLKP net1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends LARX2



.subckt LASRNX1 CLK D QN RSTB SETB VDD VSS
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net5 net3 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net3 SETB net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 QN net3 VSS VSS n12 l = 0.1u w = 0.49u m = 1
mmn3 IQN CLKP net1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net4 IQN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net6 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net5 CLKN IQN VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net1 RSTB net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmp9 QN net3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp6 net3 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 net5 RSTB VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp3 IQN CLKN net1 VDD p12 l = 0.1u w = 0.45u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp7 net5 net3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp1 net1 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net1 RSTB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net5 CLKP IQN VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 net3 IQN VDD VDD p12 l = 0.1u w = 0.39u m = 1


.ends LASRNX1



.subckt LASRNX2 CLK D QN RSTB SETB VDD VSS
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net5 net3 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net3 SETB net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 QN net3 VSS VSS n12 l = 0.1u w = 0.49u m = 2
mmn3 IQN CLKP net1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net4 IQN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net6 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net5 CLKN IQN VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net1 RSTB net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmp9 QN net3 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp6 net3 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 net5 RSTB VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp3 IQN CLKN net1 VDD p12 l = 0.1u w = 0.45u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp7 net5 net3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp1 net1 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net1 RSTB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net5 CLKP IQN VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 net3 IQN VDD VDD p12 l = 0.1u w = 0.39u m = 1


.ends LASRNX2



.subckt LASRQX1 CLK D Q RSTB SETB VDD VSS
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q net5 VSS VSS n12 l = 0.1u w = 0.49u m = 1
mmn7 net5 net3 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net3 SETB net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 IQN CLKP net1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net4 IQN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net6 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net5 CLKN IQN VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net1 RSTB net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmp6 net3 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 net5 RSTB VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp3 IQN CLKN net1 VDD p12 l = 0.1u w = 0.45u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp7 net5 net3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp1 net1 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net1 RSTB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q net5 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net5 CLKP IQN VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 net3 IQN VDD VDD p12 l = 0.1u w = 0.39u m = 1


.ends LASRQX1



.subckt LASRQX2 CLK D Q RSTB SETB VDD VSS
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q net5 VSS VSS n12 l = 0.1u w = 0.49u m = 2
mmn7 net5 net3 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net3 SETB net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 IQN CLKP net1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net4 IQN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net6 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net5 CLKN IQN VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net1 RSTB net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmp6 net3 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 net5 RSTB VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp3 IQN CLKN net1 VDD p12 l = 0.1u w = 0.45u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp7 net5 net3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp1 net1 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net1 RSTB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q net5 VDD VDD p12 l = 0.1u w = 1u m = 2
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net5 CLKP IQN VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 net3 IQN VDD VDD p12 l = 0.1u w = 0.39u m = 1


.ends LASRQX2



.subckt LASRX1 CLK D Q QN RSTB SETB VDD VSS
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q net5 VSS VSS n12 l = 0.1u w = 0.49u m = 1
mmn7 net5 net3 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net3 SETB net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 QN net3 VSS VSS n12 l = 0.1u w = 0.49u m = 1
mmn3 IQN CLKP net1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net4 IQN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net6 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net5 CLKN IQN VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net1 RSTB net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmp9 QN net3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp6 net3 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 net5 RSTB VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp3 IQN CLKN net1 VDD p12 l = 0.1u w = 0.45u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp7 net5 net3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp1 net1 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net1 RSTB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q net5 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net5 CLKP IQN VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 net3 IQN VDD VDD p12 l = 0.1u w = 0.39u m = 1


.ends LASRX1



.subckt LASRX2 CLK D Q QN RSTB SETB VDD VSS
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q net5 VSS VSS n12 l = 0.1u w = 0.56u m = 2
mmn7 net5 net3 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net3 SETB net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 QN net3 VSS VSS n12 l = 0.1u w = 0.49u m = 2
mmn3 IQN CLKP net1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net4 IQN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net6 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net5 CLKN IQN VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net1 RSTB net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmp9 QN net3 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp6 net3 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 net5 RSTB VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp3 IQN CLKN net1 VDD p12 l = 0.1u w = 0.45u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp7 net5 net3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp1 net1 D VDD VDD p12 l = 0.1u w = 0.36u m = 1
mmp2 net1 RSTB VDD VDD p12 l = 0.1u w = 0.36u m = 1
mmp10 Q net5 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net5 CLKP IQN VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 net3 IQN VDD VDD p12 l = 0.1u w = 0.39u m = 1


.ends LASRX2



.subckt LASX1 CLK D Q QN SETB VDD VSS
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 D VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q net5 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn7 net5 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net3 SETB net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 QN net3 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn3 IQN CLKP net1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net4 IQN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net5 CLKN IQN VSS n12 l = 0.1u w = 0.21u m = 1
mmp9 QN net3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp6 net3 SETB VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp7 net5 net3 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp3 IQN CLKN net1 VDD p12 l = 0.1u w = 0.4u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q net5 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net5 CLKP IQN VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 net3 IQN VDD VDD p12 l = 0.1u w = 0.35u m = 1


.ends LASX1



.subckt LASX2 CLK D Q QN SETB VDD VSS
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn1 net1 D VSS VSS n12 l = 0.1u w = 0.33u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn10 Q net5 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn7 net5 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net3 SETB net4 VSS n12 l = 0.1u w = 0.25u m = 1
mmn9 QN net3 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn3 IQN CLKP net1 VSS n12 l = 0.1u w = 0.35u m = 1
mmn5 net4 IQN VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn4 net5 CLKN IQN VSS n12 l = 0.1u w = 0.21u m = 1
mmp9 QN net3 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp6 net3 SETB VDD VDD p12 l = 0.1u w = 0.36u m = 1
mmp7 net5 net3 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp3 IQN CLKN net1 VDD p12 l = 0.1u w = 0.45u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 net1 D VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp10 Q net5 VDD VDD p12 l = 0.1u w = 2.2u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp4 net5 CLKP IQN VDD p12 l = 0.1u w = 0.21u m = 1
mmp5 net3 IQN VDD VDD p12 l = 0.1u w = 0.36u m = 1


.ends LASX2



.subckt LATCHX1 CLK D Q QN VDD VSS
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q IQN VSS VSS n12 l = 0.1u w = 0.6u m = 1
mmn7 net5 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net3 IQN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 QN net3 VSS VSS n12 l = 0.1u w = 0.6u m = 1
mmn3 IQN CLKP net1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net5 CLKN IQN VSS n12 l = 0.1u w = 0.21u m = 1
mmp9 QN net3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp5 net3 IQN VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp7 net5 net3 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp3 IQN CLKN net1 VDD p12 l = 0.1u w = 0.55u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 D VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp10 Q IQN VDD VDD p12 l = 0.1u w = 1.05u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net5 CLKP IQN VDD p12 l = 0.1u w = 0.21u m = 1


.ends LATCHX1



.subckt LATCHX2 CLK D Q QN VDD VSS
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q IQN VSS VSS n12 l = 0.1u w = 1.2u m = 1
mmn7 net5 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net3 IQN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 QN net3 VSS VSS n12 l = 0.1u w = 0.86u m = 1
mmn3 IQN CLKP net1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net5 CLKN IQN VSS n12 l = 0.1u w = 0.21u m = 1
mmp9 QN net3 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp5 net3 IQN VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp7 net5 net3 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp3 IQN CLKN net1 VDD p12 l = 0.1u w = 0.55u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 D VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp10 Q IQN VDD VDD p12 l = 0.1u w = 1.84u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net5 CLKP IQN VDD p12 l = 0.1u w = 0.21u m = 1


.ends LATCHX2



.subckt LNANDX1 Q QN RIN SIN VDD VSS
mmn3 QN Q net4 VSS n12 l = 0.1u w = 0.38u m = 1
mmn2 Q QN net2 VSS n12 l = 0.1u w = 0.38u m = 1
mmn1 net2 SIN VSS VSS n12 l = 0.1u w = 0.38u m = 1
mmn4 net4 RIN VSS VSS n12 l = 0.1u w = 0.38u m = 1
mmp2 Q QN VDD VDD p12 l = 0.1u w = 0.51u m = 1
mmp4 QN RIN VDD VDD p12 l = 0.1u w = 0.51u m = 1
mmp3 QN Q VDD VDD p12 l = 0.1u w = 0.51u m = 1
mmp1 Q SIN VDD VDD p12 l = 0.1u w = 0.51u m = 1


.ends LNANDX1



.subckt LNANDX2 Q QN RIN SIN VDD VSS
mmn3 QN Q net4 VSS n12 l = 0.1u w = 0.38u m = 2
mmn2 Q QN net2 VSS n12 l = 0.1u w = 0.38u m = 2
mmn1 net2 SIN VSS VSS n12 l = 0.1u w = 0.38u m = 2
mmn4 net4 RIN VSS VSS n12 l = 0.1u w = 0.38u m = 2
mmp2 Q QN VDD VDD p12 l = 0.1u w = 0.51u m = 2
mmp4 QN RIN VDD VDD p12 l = 0.1u w = 0.51u m = 2
mmp3 QN Q VDD VDD p12 l = 0.1u w = 0.51u m = 2
mmp1 Q SIN VDD VDD p12 l = 0.1u w = 0.51u m = 2


.ends LNANDX2



.subckt LSDNENCLSSX1 D ENB Q VDD VSS
mmn1 Q ENB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 Q ENBN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 ENBN D VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmp1 Q ENB net2 VDD p12 l = 0.1u w = 0.9u m = 1
mmp2 net2 ENBN VDD VDD p12 l = 0.1u w = 0.9u m = 1
mmp3 ENBN D VDD VDD p12 l = .1u w = .55u m = 1


.ends LSDNENCLSSX1



.subckt LSDNENCLSSX2 D ENB Q VDD VSS
mmn1 net1 D VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn2 net4 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net4 ENB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 Q net5 VSS VSS n12 l = 0.1u w = 0.56u m = 2
mmn6 net5 net4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp1 net1 D VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.9u m = 1
mmp3 net4 ENB net2 VDD p12 l = 0.1u w = 0.9u m = 1
mmp4 net5 net4 VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp6 Q net5 VDD VDD p12 l = 0.1u w = 1.1u m = 2


.ends LSDNENCLSSX2



.subckt LSDNENCLSSX4 D ENB Q VDD VSS
mmn2 111 IN2 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn1 111 ENB VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn3 IN2 D VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn6 net5 111 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 Q net5 VSS VSS n12 l = 0.1u w = 0.48u m = 4
mmp2 net2 IN2 VDD VDD p12 l = 0.1u w = 1.15u m = 1
mmp1 111 ENB net2 VDD p12 l = 0.1u w = 1.15u m = 1
mmp3 IN2 D VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp4 net5 111 VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp6 Q net5 VDD VDD p12 l = 0.1u w = 1.12u m = 4
.ends LSDNENCLSSX4



.subckt LSDNENCLSSX8 D ENB Q VDD VSS
mmn1 net1 ENB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp3 net1 VSS VSS n12 l = 0.1u w = 1.29u m = 1
mmn2 net1 ENBN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 ENBN D VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn6 Q netp3 VSS VSS n12 l = 0.1u w = 0.44u m = 8
mmp1 net1 ENB net2 VDD p12 l = 0.1u w = 0.9u m = 1
mmp2 net2 ENBN VDD VDD p12 l = 0.1u w = 0.9u m = 1
mmp3 ENBN D VDD VDD p12 l = .1u w = .55u m = 1
mmp6 netp3 net1 VDD VDD p12 l = 0.1u w = 3u m = 1
mmp7 Q netp3 VDD VDD p12 l = 0.1u w = 1.1u m = 8


.ends LSDNENCLSSX8



.subckt LSDNENCLX1 D ENB Q VDDH VDDL VSS
mmn2 Q DN VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn3 DN D VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn4 Q ENB VSS VSS n12 l = 0.1u w = 0.8u m = 1
mmp1 Q DN net2 VDDL p12 l = 0.1u w = 1.4u m = 2
mmp2 net2 ENB VDDL VDDL p12 l = 0.1u w = 1.4u m = 2
mmp3 DN D VDDH VDDH p12 l = .1u w = 0.55u m = 1


.ends LSDNENCLX1



.subckt LSDNENCLX2 D ENB Q VDDH VDDL VSS
mmp3 DN D VDDH VDDH p12 l = .1u w = 0.55u m = 1
mmp5 Q Q2 VDDL VDDL p12 l = .1u w = 3.2u m = 1
mmp2 net2 ENB VDDL VDDL p12 l = 0.1u w = 2.4u m = 1
mmp1 Q1 DN net2 VDDL p12 l = 0.1u w = 2.4u m = 1
mmp4 Q2 Q1 VDDL VDDL p12 l = .1u w = 2.8u m = 1
mmn3 DN D VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn2 Q1 DN VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn6 Q Q2 VSS VSS n12 l = 0.1u w = 1.1u m = 1
mmn5 Q2 Q1 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn4 Q1 ENB VSS VSS n12 l = 0.1u w = 0.7u m = 1


.ends LSDNENCLX2



.subckt LSDNENCLX4 D ENB Q VDDH VDDL VSS
mmp3 DN D VDDH VDDH p12 l = .1u w = 0.55u m = 1
mmp1 Q1 DN net2 VDDL p12 l = 0.1u w = 2.4u m = 1
mmp2 net2 ENB VDDL VDDL p12 l = 0.1u w = 2.4u m = 1
mmp4 Q2 Q1 VDDL VDDL p12 l = .1u w = 2.8u m = 1
mmp5 Q Q2 VDDL VDDL p12 l = .1u w = 3.2u m = 1
mmn3 DN D VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn4 Q1 ENB VSS VSS n12 l = 0.1u w = 0.7u m = 1
mmn2 Q1 DN VSS VSS n12 l = 0.1u w = 0.3u m = 1
mmn5 Q2 Q1 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn6 Q Q2 VSS VSS n12 l = 0.1u w = 1.1u m = 1


.ends LSDNENCLX4



.subckt LSDNENCLX8 D ENB Q VDDH VDDL VSS
mmp5 Q Q2 VDDL VDDL p12 l = .1u w = 3.2u m = 2
mmp2 net2 ENB VDDL VDDL p12 l = 0.1u w = 2.4u m = 1
mmp4 Q2 Q1 VDDL VDDL p12 l = .1u w = 2.8u m = 2
mmp3 DN D VDDH VDDH p12 l = .1u w = 0.55u m = 1
mmp1 Q1 DN net2 VDDL p12 l = 0.1u w = 2.4u m = 1
mmn5 Q2 Q1 VSS VSS n12 l = 0.1u w = 0.9u m = 2
mmn6 Q Q2 VSS VSS n12 l = 0.1u w = 1.1u m = 2
mmn4 Q1 ENB VSS VSS n12 l = 0.1u w = 0.7u m = 1
mmn3 DN D VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn2 Q1 DN VSS VSS n12 l = 0.1u w = 0.3u m = 1


.ends LSDNENCLX8



.subckt LSDNENSSX1 D ENB Q VDD VSS
mmn1 net1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net1 ENB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 Q net1 VSS VSS n12 l = 0.1u w = 0.48u m = 1
mmp1 net1 D net2 VDD p12 l = 0.1u w = 0.9u m = 1
mmp2 net2 ENB VDD VDD p12 l = 0.1u w = 0.9u m = 1
mmp4 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 1


.ends LSDNENSSX1



.subckt LSDNENSSX2 D ENB Q VDD VSS
mmn5 net4 net3 VSS VSS n12 l = 0.1u w = 0.48u m = 1
mmn2 net3 ENB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net3 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 Q net5 VSS VSS n12 l = 0.1u w = 0.56u m = 2
mmn6 net5 net4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 net2 ENB VDD VDD p12 l = 0.1u w = 0.9u m = 1
mmp5 net4 net3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp3 net3 D net2 VDD p12 l = 0.1u w = 0.9u m = 1
mmp4 net5 net4 VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp6 Q net5 VDD VDD p12 l = 0.1u w = 1.1u m = 2


.ends LSDNENSSX2



.subckt LSDNENSSX4 D ENB Q VDD VSS
mmn2 net1 ENB VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn5 Q net1 VSS VSS n12 l = 0.1u w = 0.48u m = 1
mmn1 net1 D VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmp2 net2 ENB VDD VDD p12 l = 0.1u w = 1.15u m = 1
mmp1 net1 D net2 VDD p12 l = 0.1u w = 1.15u m = 1
mmp5 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 1


.ends LSDNENSSX4



.subckt LSDNENSSX8 D ENB Q VDD VSS
mmn1 net1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp3 netp2 VSS VSS n12 l = 0.1u w = 1.29u m = 1
mmn2 net1 ENB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 Q netp3 VSS VSS n12 l = 0.1u w = 0.44u m = 8
mmn7 netp2 net1 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmp1 net1 D net2 VDD p12 l = 0.1u w = 0.9u m = 1
mmp2 net2 ENB VDD VDD p12 l = 0.1u w = 0.9u m = 1
mmp5 netp2 net1 VDD VDD p12 l = 0.1u w = 1u m = 1
mmp6 netp3 netp2 VDD VDD p12 l = 0.1u w = 3u m = 1
mmp7 Q netp3 VDD VDD p12 l = 0.1u w = 1.1u m = 8


.ends LSDNENSSX8



.subckt LSDNENX1 D ENB Q VDDH VDDL VSS
mmn5 net898 ENB VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn6 _n224 net898 VSS VSS n12 l = 0.1u w = 0.45u m = 1
mmn2 Q ENBN _n224 VSS n12 l = 0.1u w = 0.45u m = 1
mmn3 ENBN D VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmp1 Q ENBN VDDL VDDL p12 l = 0.1u w = 1u m = 1
mmp3 ENBN D VDDH VDDH p12 l = 0.1u w = 0.55u m = 1
mmp4 net898 ENB VDDL VDDL p12 l = 0.1u w = 0.55u m = 1
mmp5 Q net898 VDDL VDDL p12 l = 0.1u w = 1u m = 1


.ends LSDNENX1



.subckt LSDNENX2 D ENB Q VDDH VDDL VSS
mmn5 net898 ENB VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn6 _n11 net898 VSS VSS n12 l = 0.1u w = 0.44u m = 2
mmn2 Q ENBN _n11 VSS n12 l = 0.1u w = 0.44u m = 2
mmn3 ENBN D VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmp5 Q net898 VDDL VDDL p12 l = 0.1u w = 1.12u m = 2
mmp1 Q ENBN VDDL VDDL p12 l = 0.1u w = 1.12u m = 2
mmp3 ENBN D VDDH VDDH p12 l = 0.1u w = 0.55u m = 1
mmp4 net898 ENB VDDL VDDL p12 l = 0.1u w = 0.55u m = 1


.ends LSDNENX2



.subckt LSDNENX4 D ENB Q VDDH VDDL VSS
mmn6 _n76 net898 VSS VSS n12 l = 0.1u w = 0.44u m = 4
mmn2 Q ENBN _n76 VSS n12 l = 0.1u w = 0.44u m = 4
mmn3 ENBN D VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn5 net898 ENB VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmp3 ENBN D VDDH VDDH p12 l = 0.1u w = 0.55u m = 1
mmp5 Q net898 VDDL VDDL p12 l = 0.1u w = 1u m = 4
mmp1 Q ENBN VDDL VDDL p12 l = 0.1u w = 1u m = 4
mmp4 net898 ENB VDDL VDDL p12 l = 0.1u w = 0.55u m = 1


.ends LSDNENX4



.subckt LSDNENX8 D ENB Q VDDH VDDL VSS


mmp3 ENBN D VDDH VDDH p12 l = 0.1u w = 0.55u m = 1
mmp1 Q ENBN VDDL VDDL p12 l = 0.1u w = 1.12u m = 8
mmp4 net898 ENB VDDL VDDL p12 l = 0.1u w = 0.55u m = 1
mmp5 Q net898 VDDL VDDL p12 l = 0.1u w = 1.12u m = 8
mmn2 Q ENBN _n173 VSS n12 l = 0.1u w = 0.44u m = 8
mmn6 _n173 net898 VSS VSS n12 l = 0.1u w = 0.44u m = 8
mmn3 ENBN D VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn5 net898 ENB VSS VSS n12 l = 0.1u w = 0.24u m = 1
.ends LSDNENX8



.subckt LSDNSSX1 D Q VDD VSS
mmn2 Q netp1 VSS VSS n12 l = 0.1u w = 0.49u m = 1
mmn1 netp1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 Q netp1 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp1 netp1 D VDD VDD p12 l = 0.1u w = 0.5u m = 1


.ends LSDNSSX1



.subckt LSDNSSX2 D Q VDD VSS
mmn2 Q netp1 VSS VSS n12 l = 0.1u w = 0.56u m = 2
mmn1 netp1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 Q netp1 VDD VDD p12 l = 0.1u w = 1.1u m = 2
mmp1 netp1 D VDD VDD p12 l = 0.1u w = 0.55u m = 1


.ends LSDNSSX2



.subckt LSDNSSX4 D Q VDD VSS
mmn2 Q netp1 VSS VSS n12 l = 0.1u w = 0.475u m = 4
mmn1 netp1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 Q netp1 VDD VDD p12 l = 0.1u w = 1.05u m = 4
mmp1 netp1 D VDD VDD p12 l = 0.1u w = 0.6u m = 1


.ends LSDNSSX4



.subckt LSDNSSX8 D Q VDD VSS
mmn2 netp2 netp1 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn1 netp1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 netp3 netp2 VSS VSS n12 l = 0.1u w = 1.29u m = 1
mmn4 Q netp3 VSS VSS n12 l = 0.1u w = 0.44u m = 8
mmp2 netp2 netp1 VDD VDD p12 l = 0.1u w = 1u m = 1
mmp1 netp1 D VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp3 netp3 netp2 VDD VDD p12 l = 0.1u w = 3u m = 1
mmp4 Q netp3 VDD VDD p12 l = 0.1u w = 1.1u m = 8


.ends LSDNSSX8



.subckt LSDNX1 D Q VDDH VDDL VSS
mmn2 Q netp1 VSS VSS n12 l = 0.1u w = 0.49u m = 1
mmn1 netp1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 Q netp1 VDDL VDDL p12 l = 0.1u w = 1.12u m = 1
mmp1 netp1 D VDDH VDDH p12 l = 0.1u w = 0.5u m = 1


.ends LSDNX1



.subckt LSDNX2 D Q VDDH VDDL VSS
mmn2 Q netp1 VSS VSS n12 l = 0.1u w = 0.56u m = 2
mmn1 netp1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 Q netp1 VDDL VDDL p12 l = 0.1u w = 1.1u m = 2
mmp1 netp1 D VDDH VDDH p12 l = 0.1u w = 0.55u m = 1


.ends LSDNX2



.subckt LSDNX4 D Q VDDH VDDL VSS
mmn2 Q netp1 VSS VSS n12 l = 0.1u w = 0.475u m = 4
mmn1 netp1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 Q netp1 VDDL VDDL p12 l = 0.1u w = 1.05u m = 4
mmp1 netp1 D VDDH VDDH p12 l = 0.1u w = 0.6u m = 1


.ends LSDNX4



.subckt LSDNX8 D Q VDDH VDDL VSS


mmp1 netp1 D VDDH VDDH p12 l = 0.1u w = 0.21u m = 1
mmp2 netp2 netp1 VDDL VDDL p12 l = 0.1u w = 1u m = 1
mmp3 netp3 netp2 VDDL VDDL p12 l = 0.1u w = 3u m = 1
mmp4 Q netp3 VDDL VDDL p12 l = 0.1u w = 1.1u m = 8
mmn1 netp1 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netp2 netp1 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn3 netp3 netp2 VSS VSS n12 l = 0.1u w = 1.29u m = 1
mmn4 Q netp3 VSS VSS n12 l = 0.1u w = 0.44u m = 8
.ends LSDNX8



.subckt LSUPENCLX1 D ENB Q VDDH VDDL VSS
mmp1 net1 D VDDL VDDL p12 l = 0.1u w = 0.22u m = 1
mmp3 net4 net3 mm VDDH p12 l = 0.1u w = 0.5u m = 1
mmp4 Q net4 mm VDDH p12 l = 0.1u w = 1.12u m = 1
mmp2 net3 net4 mm VDDH p12 l = 0.1u w = 0.5u m = 1
mmp5 mm ENB VDDH VDDH p12 l = 0.1u w = 0.8u m = 1
mmn1 net1 D VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn3 net4 D VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn4 Q net4 VSS VSS n12 l = 0.1u w = 0.55u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.28u m = 1
mmn6 Q ENB VSS VSS n12 l = 0.1u w = 0.8u m = 1


.ends LSUPENCLX1



.subckt LSUPENCLX2 D ENB Q VDDH VDDL VSS
mmp4 Q net3 _n34 VDDH p12 l = 0.1u w = 1u m = 2
mmp2 net2 net3 _n34 VDDH p12 l = 0.1u w = 0.54u m = 1
mmp1 net1 D VDDL VDDL p12 l = 0.1u w = 0.22u m = 1
mmp3 net3 net2 _n34 VDDH p12 l = 0.1u w = 0.54u m = 1
mmp5 _n34 ENB VDDH VDDH p12 l = 0.1u w = 1u m = 1
mmn4 Q net3 VSS VSS n12 l = 0.1u w = 0.35u m = 2
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.28u m = 1
mmn3 net3 D VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn1 net1 D VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn5 Q ENB VSS VSS n12 l = 0.1u w = 0.4u m = 1


.ends LSUPENCLX2



.subckt LSUPENCLX4 D ENB Q VDDH VDDL VSS
mmp1 net1 D VDDL VDDL p12 l = 0.1u w = 0.22u m = 1
mmp3 net4 net3 _n29 VDDH p12 l = 0.1u w = 0.5u m = 1
mmp4 Q net4 _n29 VDDH p12 l = 0.1u w = 1.4u m = 4
mmp2 net3 net4 _n29 VDDH p12 l = 0.1u w = 0.5u m = 1
mmp5 _n29 ENB VDDH VDDH p12 l = 0.1u w = 0.8u m = 1
mmn1 net1 D VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn3 net4 D VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn4 Q net4 VSS VSS n12 l = 0.1u w = 1.1u m = 4
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.28u m = 1
mmn6 Q ENB VSS VSS n12 l = 0.1u w = 0.8u m = 1


.ends LSUPENCLX4



.subckt LSUPENCLX8 D ENB Q VDDH VDDL VSS
mmp1 net1 D VDDL VDDL p12 l = 0.1u w = 0.22u m = 1
mmp3 net4 net3 _n29 VDDH p12 l = 0.1u w = 0.5u m = 1
mmp4 Q net4 _n29 VDDH p12 l = 0.1u w = 2.4u m = 8
mmp2 net3 net4 _n29 VDDH p12 l = 0.1u w = 0.5u m = 1
mmp5 _n29 ENB VDDH VDDH p12 l = 0.1u w = 3.5u m = 1
mmn1 net1 D VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn3 net4 D VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn4 Q net4 VSS VSS n12 l = 0.1u w = 1.6u m = 8
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.7u m = 1
mmn6 Q ENB VSS VSS n12 l = 0.1u w = 2.5u m = 1


.ends LSUPENCLX8



.subckt LSUPENX1 D ENB Q VDDH VDDL VSS
mmp1 net1 D VDDL VDDL p12 l = 0.1u w = 0.22u m = 1
mmp3 net4 net3 VDDH VDDH p12 l = 0.1u w = 0.4u m = 1
mmp4 Q net4 VDDH VDDH p12 l = 0.1u w = 0.54u m = 1
mmp2 net3 net4 VDDH VDDH p12 l = 0.1u w = 0.4u m = 1
mmp5 Q net98 VDDH VDDH p12 l = 0.1u w = 0.8u m = 2
mmp6 net98 ENB VDDH VDDH p12 l = 0.1u w = 0.22u m = 1
mmn1 net1 D VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn3 net4 D net2 VSS n12 l = 0.1u w = 0.25u m = 1
mmn4 Q net4 net2 VSS n12 l = 0.1u w = 0.23u m = 1
mmn2 net3 net1 net2 VSS n12 l = 0.1u w = 0.25u m = 1
mmn5 net2 net98 VSS VSS n12 l = 0.1u w = 0.8u m = 2
mmn6 net98 ENB VSS VSS n12 l = 0.1u w = 0.22u m = 1


.ends LSUPENX1



.subckt LSUPENX2 D ENB Q VDDH VDDL VSS
mmp4 Q net3 VDDH VDDH p12 l = 0.1u w = 0.4u m = 2
mmp2 net2 net3 VDDH VDDH p12 l = 0.1u w = 0.36u m = 1
mmp1 net1236 D VDDL VDDL p12 l = 0.1u w = 0.22u m = 1
mmp3 net3 net2 VDDH VDDH p12 l = 0.1u w = 0.36u m = 1
mmp5 net1 ENB VDDH VDDH p12 l = 0.1u w = 0.22u m = 1
mmp6 Q net1 VDDH VDDH p12 l = 0.1u w = 2.24u m = 1
mmn4 Q net3 net4 VSS n12 l = 0.1u w = 0.2u m = 2
mmn2 net2 net1236 net4 VSS n12 l = 0.1u w = 0.28u m = 1
mmn3 net3 D net4 VSS n12 l = 0.1u w = 0.25u m = 1
mmn1 net1236 D VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn5 net4 net1 VSS VSS n12 l = 0.1u w = 2.24u m = 1
mmn6 net1 ENB VSS VSS n12 l = 0.1u w = 0.22u m = 1


.ends LSUPENX2



.subckt LSUPENX4 D ENB Q VDDH VDDL VSS
mmp5 Q net98 VDDH VDDH p12 l = 0.1u w = 1.1u m = 2
mmp4 Q net3 VDDH VDDH p12 l = 0.1u w = 1.12u m = 4
mmp3 net3 net2 VDDH VDDH p12 l = 0.1u w = 0.61u m = 1
mmp2 VDDH net3 net2 VDDH p12 l = 0.1u w = 0.61u m = 1
mmp1 net1 D VDDL VDDL p12 l = 0.1u w = 0.46u m = 1
mmp6 net98 ENB VDDH VDDH p12 l = 0.1u w = 0.46u m = 1
mmn1 net1 D VSS VSS n12 l = 0.1u w = 0.46u m = 1
mmn3 net3 D net0 VSS n12 l = 0.1u w = 0.51u m = 1
mmn2 net2 net1 net0 VSS n12 l = 0.1u w = 0.51u m = 1
mmn4 Q net3 net0 VSS n12 l = 0.1u w = 0.64u m = 4
mmn5 net0 net98 VSS VSS n12 l = 0.1u w = 1.1u m = 2
mmn6 net98 ENB VSS VSS n12 l = 0.1u w = 0.46u m = 1
.ends LSUPENX4



.subckt LSUPENX8 D ENB Q VDDH VDDL VSS


mmp4 Q net3 VDDH VDDH p12 l = 0.1u w = 1.12u m = 8
mmp1 net1 D VDDL VDDL p12 l = 0.1u w = 0.46u m = 1
mmp2 VDDH net3 net2 VDDH p12 l = 0.1u w = 0.455u m = 1
mmp3 net3 net2 VDDH VDDH p12 l = 0.1u w = 0.455u m = 1
mmp5 Q netp VDDH VDDH p12 l = 0.1u w = 1.1u m = 2
mmp6 netp ENB VDDH VDDH p12 l = 0.1u w = 0.46u m = 1
mmn1 net1 D VSS VSS n12 l = 0.1u w = 0.46u m = 1
mmn5 net0 netp VSS VSS n12 l = 0.1u w = 1.1u m = 2
mmn4 Q net3 net0 VSS n12 l = 0.1u w = 0.62u m = 8
mmn2 net2 net1 net0 VSS n12 l = 0.1u w = 0.41u m = 1
mmn3 net3 D net0 VSS n12 l = 0.1u w = 0.41u m = 1
mmn6 netp ENB VSS VSS n12 l = 0.1u w = 0.46u m = 1
.ends LSUPENX8



.subckt LSUPX1 D Q VDDH VDDL VSS
mmp1 mp1 D VDDL VDDL p12 l = 0.1u w = 0.22u m = 1
mmp3 mp3 mp2 VDDH VDDH p12 l = 0.1u w = 0.4u m = 1
mmp4 Q mp3 VDDH VDDH p12 l = 0.1u w = 1.12u m = 1
mmp2 mp2 mp3 VDDH VDDH p12 l = 0.1u w = 0.4u m = 1
mmn1 mp1 D VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn3 mp3 D VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn4 Q mp3 VSS VSS n12 l = 0.1u w = 0.55u m = 1
mmn2 mp2 mp1 VSS VSS n12 l = 0.1u w = 0.25u m = 1


.ends LSUPX1



.subckt LSUPX2 D Q VDDH VDDL VSS
mmp1 mp1 D VDDL VDDL p12 l = 0.1u w = 0.22u m = 1
mmp3 mp3 mp2 VDDH VDDH p12 l = 0.1u w = 0.4u m = 1
mmp4 Q mp3 VDDH VDDH p12 l = 0.1u w = 1.12u m = 2
mmp2 mp2 mp3 VDDH VDDH p12 l = 0.1u w = 0.4u m = 1
mmn1 mp1 D VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn3 mp3 D VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn4 Q mp3 VSS VSS n12 l = 0.1u w = 0.55u m = 2
mmn2 mp2 mp1 VSS VSS n12 l = 0.1u w = 0.25u m = 1


.ends LSUPX2



.subckt LSUPX4 D Q VDDH VDDL VSS
mmp1 mp1 D VDDL VDDL p12 l = 0.1u w = 0.22u m = 1
mmp3 mp3 mp2 VDDH VDDH p12 l = 0.1u w = 0.4u m = 1
mmp4 Q mp3 VDDH VDDH p12 l = 0.1u w = 1.12u m = 4
mmp2 mp2 mp3 VDDH VDDH p12 l = 0.1u w = 0.4u m = 1
mmn1 mp1 D VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn3 mp3 D VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn4 Q mp3 VSS VSS n12 l = 0.1u w = 0.55u m = 4
mmn2 mp2 mp1 VSS VSS n12 l = 0.1u w = 0.25u m = 1


.ends LSUPX4



.subckt LSUPX8 D Q VDDH VDDL VSS
mmp1 mp1 D VDDL VDDL p12 l = 0.1u w = 0.22u m = 1
mmp3 mp3 mp2 VDDH VDDH p12 l = 0.1u w = 0.4u m = 1
mmp4 Q mp3 VDDH VDDH p12 l = 0.1u w = 1.12u m = 8
mmp2 mp2 mp3 VDDH VDDH p12 l = 0.1u w = 0.4u m = 1
mmn1 mp1 D VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn3 mp3 D VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn4 Q mp3 VSS VSS n12 l = 0.1u w = 0.55u m = 8
mmn2 mp2 mp1 VSS VSS n12 l = 0.1u w = 0.25u m = 1


.ends LSUPX8



.subckt MUX21X1 IN1 IN2 Q S VDD VSS
mmp1 net1 S VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp5 net3 IN2 net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmp4 net5 net1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp3 net3 IN1 net2 VDD p12 l = 0.1u w = 0.65u m = 1
mmp6 Q net3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp2 net2 S VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmn3 net4 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 IN1 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 S VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net6 S VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 Q net3 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn4 net3 IN2 net6 VSS n12 l = 0.1u w = 0.21u m = 1


.ends MUX21X1



.subckt MUX21X2 IN1 IN2 Q S VDD VSS
mmp1 net1 S VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp5 net3 IN2 net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmp4 net5 net1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp3 net3 IN1 net2 VDD p12 l = 0.1u w = 0.65u m = 1
mmp6 Q net3 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp2 net2 S VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmn3 net4 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 IN1 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 S VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net6 S VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 Q net3 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn4 net3 IN2 net6 VSS n12 l = 0.1u w = 0.21u m = 1


.ends MUX21X2



.subckt MUX41X1 IN1 IN2 IN3 IN4 Q S0 S1 VDD VSS
mmp1 net1 S1 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp2 net4 IN1 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp3 net2 S1 net4 VDD p12 l = 0.1u w = 0.6u m = 1
mmp4 net6 IN2 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp5 net2 net1 net6 VDD p12 l = 0.1u w = 0.6u m = 1
mmp6 net3 S1 net10 VDD p12 l = 0.1u w = 0.6u m = 1
mmp7 net10 IN3 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp8 net3 net1 net12 VDD p12 l = 0.1u w = 0.6u m = 1
mmp9 net12 IN4 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp10 net7 S0 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp11 net2 S0 net8 VDD p12 l = 0.1u w = 0.55u m = 1
mmp12 net3 net7 net8 VDD p12 l = 0.1u w = 0.55u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmn1 net1 S1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net5 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net2 S1 net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net9 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net3 net1 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net11 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net3 S1 net13 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net13 IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net7 S0 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net2 net7 net8 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net3 S0 net8 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.43u m = 1


.ends MUX41X1



.subckt MUX41X2 IN1 IN2 IN3 IN4 Q S0 S1 VDD VSS
mmp1 net1 S1 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp2 net4 IN1 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp3 net2 S1 net4 VDD p12 l = 0.1u w = 0.6u m = 1
mmp4 net6 IN2 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp5 net2 net1 net6 VDD p12 l = 0.1u w = 0.6u m = 1
mmp6 net3 S1 net10 VDD p12 l = 0.1u w = 0.6u m = 1
mmp7 net10 IN3 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp8 net3 net1 net12 VDD p12 l = 0.1u w = 0.6u m = 1
mmp9 net12 IN4 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp10 net7 S0 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp11 net2 S0 net8 VDD p12 l = 0.1u w = 0.7u m = 1
mmp12 net3 net7 net8 VDD p12 l = 0.1u w = 0.7u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmn1 net1 S1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net5 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net2 S1 net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net9 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net3 net1 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net11 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net3 S1 net13 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net13 IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net7 S0 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net2 net7 net8 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net3 S0 net8 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.43u m = 2


.ends MUX41X2



.subckt NAND2X0 IN1 IN2 QN VDD VSS
mmp3 QN IN2 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp4 QN IN1 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmn3 net1 IN2 VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn4 QN IN1 net1 VSS n12 l = 0.1u w = 0.25u m = 1


.ends NAND2X0



.subckt NAND2X1 IN1 IN2 QN VDD VSS
mmn2 net1 IN2 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn1 QN IN1 net1 VSS n12 l = 0.1u w = 0.5u m = 1
mmp2 QN IN2 VDD VDD p12 l = 0.1u w = 0.8u m = 1
mmp1 QN IN1 VDD VDD p12 l = 0.1u w = 0.8u m = 1


.ends NAND2X1



.subckt NAND2X2 IN1 IN2 QN VDD VSS
mmn3 net1 IN2 VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn4 QN IN1 net1 VSS n12 l = 0.1u w = 0.5u m = 2
mmp3 QN IN2 VDD VDD p12 l = 0.1u w = 0.8u m = 2
mmp4 QN IN1 VDD VDD p12 l = 0.1u w = 0.8u m = 2


.ends NAND2X2



.subckt NAND2X4 IN1 IN2 QN VDD VSS
mmn3 net1 IN2 VSS VSS n12 l = 0.1u w = 0.5u m = 4
mmn4 QN IN1 net1 VSS n12 l = 0.1u w = 0.5u m = 4
mmp3 QN IN2 VDD VDD p12 l = 0.1u w = 0.8u m = 4
mmp4 QN IN1 VDD VDD p12 l = 0.1u w = 0.8u m = 4


.ends NAND2X4



.subckt NAND3X0 IN1 IN2 IN3 QN VDD VSS
mmn2 net1 IN2 net2 VSS n12 l = 0.1u w = 0.52u m = 1
mmn3 net2 IN3 VSS VSS n12 l = 0.1u w = 0.52u m = 1
mmn1 QN IN1 net1 VSS n12 l = 0.1u w = 0.52u m = 1
mmp1 QN IN1 VDD VDD p12 l = 0.1u w = 0.58u m = 1
mmp2 QN IN2 VDD VDD p12 l = 0.1u w = 0.58u m = 1
mmp3 QN IN3 VDD VDD p12 l = 0.1u w = 0.58u m = 1


.ends NAND3X0



.subckt NAND3X1 IN1 IN2 IN3 QN VDD VSS
mmn2 net1 IN2 net2 VSS n12 l = 0.1u w = 0.28u m = 1
mmn1 net4 IN1 net1 VSS n12 l = 0.1u w = 0.28u m = 1
mmn3 net2 IN3 VSS VSS n12 l = 0.1u w = 0.28u m = 1
mmn4 net5 net4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 QN net5 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmp2 net4 IN2 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp3 net4 IN3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp4 net5 net4 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp1 net4 IN1 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp5 QN net5 VDD VDD p12 l = 0.1u w = 1.12u m = 1


.ends NAND3X1



.subckt NAND3X2 IN1 IN2 IN3 QN VDD VSS
mmp6 QN net5 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp7 net4 IN3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp8 net4 IN1 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp9 net4 IN2 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp10 net5 net4 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmn6 net4 IN1 net1 VSS n12 l = 0.1u w = 0.28u m = 1
mmn7 QN net5 VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn8 net1 IN2 net2 VSS n12 l = 0.1u w = 0.28u m = 1
mmn9 net2 IN3 VSS VSS n12 l = 0.1u w = 0.28u m = 1
mmn10 net5 net4 VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends NAND3X2



.subckt NAND3X4 IN1 IN2 IN3 QN VDD VSS
mmp6 QN net5 VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmp7 net4 IN3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp8 net4 IN1 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp9 net4 IN2 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp10 net5 net4 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmn6 net4 IN1 net1 VSS n12 l = 0.1u w = 0.28u m = 1
mmn7 QN net5 VSS VSS n12 l = 0.1u w = 0.5u m = 4
mmn8 net1 IN2 net2 VSS n12 l = 0.1u w = 0.28u m = 1
mmn9 net2 IN3 VSS VSS n12 l = 0.1u w = 0.28u m = 1
mmn10 net5 net4 VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends NAND3X4



.subckt NAND4X0 IN1 IN2 IN3 IN4 QN VDD VSS
mmn3 net2 IN3 net3 VSS n12 l = 0.1u w = 0.53u m = 1
mmn1 QN IN1 net1 VSS n12 l = 0.1u w = 0.53u m = 1
mmn4 net3 IN4 VSS VSS n12 l = 0.1u w = 0.53u m = 1
mmn2 net1 IN2 net2 VSS n12 l = 0.1u w = 0.53u m = 1
mmp1 QN IN1 VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp2 QN IN2 VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp4 QN IN4 VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 QN IN3 VDD VDD p12 l = 0.1u w = 0.48u m = 1


.ends NAND4X0



.subckt NAND4X1 IN1 IN2 IN3 IN4 QN VDD VSS
mmp2 net1 IN2 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp3 net1 IN3 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp4 net1 IN4 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp5 net5 net1 VDD VDD p12 l = 0.1u w = 0.63u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp6 QN net5 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmn1 net1 IN1 net2 VSS n12 l = 0.1u w = 0.5u m = 1
mmn2 net2 IN2 net3 VSS n12 l = 0.1u w = 0.5u m = 1
mmn3 net3 IN3 net4 VSS n12 l = 0.1u w = 0.5u m = 1
mmn4 net4 IN4 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn5 net5 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 QN net5 VSS VSS n12 l = 0.1u w = 0.4u m = 1


.ends NAND4X1



.subckt NBUFFX16 INP VDD VSS Z
mmp2 Z net1 VDD VDD p12 l = 0.1u w = 1.12u m = 16
mmp1 net1 INP VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmn1 net1 INP VSS VSS n12 l = 0.1u w = 0.37u m = 2
mmn2 Z net1 VSS VSS n12 l = 0.1u w = 0.43u m = 16


.ends NBUFFX16



.subckt NBUFFX2 INP VDD VSS Z
mmn2 Z net1 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn1 net1 INP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 Z net1 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp1 net1 INP VDD VDD p12 l = 0.1u w = 0.62u m = 1


.ends NBUFFX2



.subckt NBUFFX32 INP VDD VSS Z
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp1 net1 INP VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp4 Z net3 VDD VDD p12 l = 0.1u w = 1.12u m = 32
mmp3 net3 net2 VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmn1 net1 INP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn4 Z net3 VSS VSS n12 l = 0.1u w = 0.43u m = 32
mmn3 net3 net2 VSS VSS n12 l = 0.1u w = 0.43u m = 4


.ends NBUFFX32



.subckt NBUFFX4 INP VDD VSS Z
mmp2 Z net1 VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmp1 net1 INP VDD VDD p12 l = 0.1u w = 0.62u m = 1
mmn2 Z net1 VSS VSS n12 l = 0.1u w = 0.43u m = 4
mmn1 net1 INP VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends NBUFFX4



.subckt NBUFFX8 INP VDD VSS Z
mmp1 net1 INP VDD VDD p12 l = 0.1u w = 1.17u m = 1
mmp2 Z net1 VDD VDD p12 l = 0.1u w = 1.12u m = 8
mmn1 net1 INP VSS VSS n12 l = 0.1u w = 0.38u m = 1
mmn2 Z net1 VSS VSS n12 l = 0.1u w = 0.43u m = 8


.ends NBUFFX8



.subckt NMT1 D G S VDD VSS


mg_nmos4t1 D G S VSS n12 l = 0.1u w = 0.48u m = 1
.ends NMT1



.subckt NMT2 D G S VDD VSS


mg_nmos4t1 D G S VSS n12 l = 0.1u w = 0.48u m = 2
.ends NMT2



.subckt NMT3 D G S VDD VSS
mg_nmos4t1 D G S VSS n12 l = 0.1u w = 0.48u m = 4


.ends NMT3



.subckt NOR2X0 IN1 IN2 QN VDD VSS
mmp3 net2 IN2 VDD VDD p12 l = 0.1u w = 0.8u m = 1
mmp4 QN IN1 net2 VDD p12 l = 0.1u w = 0.8u m = 1
mmn3 QN IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 QN IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends NOR2X0



.subckt NOR2X1 IN1 IN2 QN VDD VSS
mmn1 QN IN1 VSS VSS n12 l = 0.1u w = 0.28u m = 1
mmn2 QN IN2 VSS VSS n12 l = 0.1u w = 0.28u m = 1
mmp2 net2 IN2 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp1 QN IN1 net2 VDD p12 l = 0.1u w = 1.12u m = 1


.ends NOR2X1



.subckt NOR2X2 IN1 IN2 QN VDD VSS
mmp3 net2 IN2 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp4 QN IN1 net2 VDD p12 l = 0.1u w = 1.12u m = 2
mmn3 QN IN1 VSS VSS n12 l = 0.1u w = 0.28u m = 2
mmn4 QN IN2 VSS VSS n12 l = 0.1u w = 0.28u m = 2


.ends NOR2X2



.subckt NOR2X4 IN1 IN2 QN VDD VSS
mmn3 QN IN1 VSS VSS n12 l = 0.1u w = 0.28u m = 4
mmn4 QN IN2 VSS VSS n12 l = 0.1u w = 0.28u m = 4
mmp3 net2 IN2 VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmp4 QN IN1 net2 VDD p12 l = 0.1u w = 1.12u m = 4


.ends NOR2X4



.subckt NOR3X0 IN1 IN2 IN3 QN VDD VSS
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp1 QN IN1 net2 VDD p12 l = 0.1u w = 1.12u m = 1
mmp2 net2 IN2 net3 VDD p12 l = 0.1u w = 1.12u m = 1
mmn3 QN IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 QN IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 QN IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends NOR3X0



.subckt NOR3X1 IN1 IN2 IN3 QN VDD VSS
mmn2 net1 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net1 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net5 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 QN net5 VSS VSS n12 l = 0.1u w = 0.54u m = 1
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp1 net1 IN1 net2 VDD p12 l = 0.1u w = 1.12u m = 1
mmp2 net2 IN2 net3 VDD p12 l = 0.1u w = 1.12u m = 1
mmp4 net5 net1 VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp5 QN net5 VDD VDD p12 l = 0.1u w = 1.12u m = 1


.ends NOR3X1



.subckt NOR3X2 IN1 IN2 IN3 QN VDD VSS
mmn6 net1 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net1 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net5 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net1 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 QN net5 VSS VSS n12 l = 0.1u w = 0.54u m = 2
mmp6 net2 IN2 net3 VDD p12 l = 0.1u w = 1.12u m = 1
mmp7 net5 net1 VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp8 net3 IN3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp9 QN net5 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp10 net1 IN1 net2 VDD p12 l = 0.1u w = 1.12u m = 1


.ends NOR3X2



.subckt NOR3X4 IN1 IN2 IN3 QN VDD VSS
mmn7 net1 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 QN net5 VSS VSS n12 l = 0.1u w = 0.54u m = 4
mmn8 net5 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net1 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp7 net5 net1 VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp10 net1 IN1 net2 VDD p12 l = 0.1u w = 1.12u m = 1
mmp8 net3 IN3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp6 net2 IN2 net3 VDD p12 l = 0.1u w = 1.12u m = 1
mmp9 QN net5 VDD VDD p12 l = 0.1u w = 1.12u m = 4


.ends NOR3X4



.subckt NOR4X0 IN1 IN2 IN3 IN4 QN VDD VSS
mmp3 net3 IN3 net4 VDD p12 l = 0.1u w = 1.12u m = 1
mmp2 net2 IN2 net3 VDD p12 l = 0.1u w = 1.12u m = 1
mmp4 net4 IN4 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp1 QN IN1 net2 VDD p12 l = 0.1u w = 1.12u m = 1
mmn1 QN IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 QN IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 QN IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 QN IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends NOR4X0



.subckt NOR4X1 IN1 IN2 IN3 IN4 QN VDD VSS
mmn2 net3 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net3 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net4 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net4 IN4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net6 net3 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net5 net4 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 QN net6 VSS VSS n12 l = 0.1u w = 0.45u m = 1
mmp2 net1 IN1 VDD VDD p12 l = 0.1u w = 0.75u m = 1
mmp1 net3 IN2 net1 VDD p12 l = 0.1u w = 0.75u m = 1
mmp3 net2 IN3 VDD VDD p12 l = 0.1u w = 0.75u m = 1
mmp4 net4 IN4 net2 VDD p12 l = 0.1u w = 0.75u m = 1
mmp5 net6 net4 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp6 net6 net3 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp7 QN net6 VDD VDD p12 l = 0.1u w = 1.12u m = 1


.ends NOR4X1



.subckt OA21X1 IN1 IN2 IN3 Q VDD VSS
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn4 Q net3 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn3 net3 IN3 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp4 Q net3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp2 net3 IN2 net1 VDD p12 l = 0.1u w = 0.55u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.55u m = 1


.ends OA21X1



.subckt OA21X2 IN1 IN2 IN3 Q VDD VSS
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp2 net3 IN2 net1 VDD p12 l = 0.1u w = 0.68u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.68u m = 1
mmp4 Q net3 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmn4 Q net3 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net3 IN3 net2 VSS n12 l = 0.1u w = 0.21u m = 1


.ends OA21X2



.subckt OA221X1 IN1 IN2 IN3 IN4 IN5 Q VDD VSS
mmp6 Q net5 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp5 net5 IN5 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.58u m = 1
mmp2 net5 IN2 net1 VDD p12 l = 0.1u w = 0.58u m = 1
mmp4 net5 IN4 net3 VDD p12 l = 0.1u w = 0.55u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net4 IN4 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net4 IN3 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 Q net5 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn5 net5 IN5 net4 VSS n12 l = 0.1u w = 0.3u m = 1


.ends OA221X1



.subckt OA221X2 IN1 IN2 IN3 IN4 IN5 Q VDD VSS
mmp5 net5 IN5 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp4 net5 IN4 net3 VDD p12 l = 0.1u w = 0.55u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.57u m = 1
mmp6 Q net5 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp2 net5 IN2 net1 VDD p12 l = 0.1u w = 0.57u m = 1
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmn4 net4 IN4 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 IN5 net4 VSS n12 l = 0.1u w = 0.3u m = 1
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 Q net5 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn3 net4 IN3 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends OA221X2



.subckt OA222X1 IN1 IN2 IN3 IN4 IN5 IN6 Q VDD VSS
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net4 IN3 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net6 IN6 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net6 IN5 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net4 IN4 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 Q net6 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.45u m = 1
mmp5 net5 IN5 VDD VDD p12 l = 0.1u w = 0.45u m = 1
mmp6 net6 IN6 net5 VDD p12 l = 0.1u w = 0.45u m = 1
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.45u m = 1
mmp4 net6 IN4 net3 VDD p12 l = 0.1u w = 0.45u m = 1
mmp2 net6 IN2 net1 VDD p12 l = 0.1u w = 0.6u m = 1
mmp7 Q net6 VDD VDD p12 l = 0.1u w = 1.12u m = 1


.ends OA222X1



.subckt OA222X2 IN1 IN2 IN3 IN4 IN5 IN6 Q VDD VSS
mmp2 net6 IN2 net1 VDD p12 l = 0.1u w = 0.6u m = 1
mmp5 net5 IN5 VDD VDD p12 l = 0.1u w = 0.45u m = 1
mmp4 net6 IN4 net3 VDD p12 l = 0.1u w = 0.45u m = 1
mmp7 Q net6 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp6 net6 IN6 net5 VDD p12 l = 0.1u w = 0.45u m = 1
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.45u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.45u m = 1
mmn3 net4 IN3 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net6 IN5 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net6 IN6 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net4 IN4 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 Q net6 VSS VSS n12 l = 0.1u w = 0.43u m = 2


.ends OA222X2



.subckt OA22X1 IN1 IN2 IN3 IN4 Q VDD VSS
mmn5 Q net4 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn4 net4 IN4 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net4 IN3 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp4 net4 IN4 net3 VDD p12 l = 0.1u w = 0.58u m = 1
mmp5 Q net4 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.7u m = 1
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.58u m = 1
mmp2 net4 IN2 net1 VDD p12 l = 0.1u w = 0.7u m = 1


.ends OA22X1



.subckt OA22X2 IN1 IN2 IN3 IN4 Q VDD VSS
mmn3 net4 IN3 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net4 IN4 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 Q net4 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp4 net4 IN4 net3 VDD p12 l = 0.1u w = 0.58u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.7u m = 1
mmp5 Q net4 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.58u m = 1
mmp2 net4 IN2 net1 VDD p12 l = 0.1u w = 0.7u m = 1


.ends OA22X2



.subckt OAI21X1 IN1 IN2 IN3 QN VDD VSS
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn4 net4 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net3 IN3 net2 VSS n12 l = 0.1u w = 0.32u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn5 QN net4 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net3 IN2 net1 VDD p12 l = 0.1u w = 0.48u m = 1
mmp4 net4 net3 VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp5 QN net4 VDD VDD p12 l = 0.1u w = 1.12u m = 1


.ends OAI21X1



.subckt OAI21X2 IN1 IN2 IN3 QN VDD VSS
mmn5 QN net4 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn3 net3 IN3 net2 VSS n12 l = 0.1u w = 0.32u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn4 net4 net3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp5 QN net4 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp2 net3 IN2 net1 VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net4 net3 VDD VDD p12 l = 0.1u w = 0.55u m = 1


.ends OAI21X2



.subckt OAI221X1 IN1 IN2 IN3 IN4 IN5 QN VDD VSS
mmp7 QN net6 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp2 net5 IN2 net1 VDD p12 l = 0.1u w = 0.4u m = 1
mmp5 net5 IN5 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net5 IN4 net3 VDD p12 l = 0.1u w = 0.4u m = 1
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp6 net6 net5 VDD VDD p12 l = 0.1u w = 0.37u m = 1
mmn7 QN net6 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn4 net4 IN4 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn3 net4 IN3 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn6 net6 net5 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn5 net5 IN5 net4 VSS n12 l = 0.1u w = 0.25u m = 1


.ends OAI221X1



.subckt OAI221X2 IN1 IN2 IN3 IN4 IN5 QN VDD VSS
mmn5 net5 IN5 net4 VSS n12 l = 0.1u w = 0.25u m = 1
mmn6 net6 net5 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn4 net4 IN4 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 QN net6 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn3 net4 IN3 net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmp6 net6 net5 VDD VDD p12 l = 0.1u w = 0.37u m = 1
mmp7 QN net6 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp2 net5 IN2 net1 VDD p12 l = 0.1u w = 0.4u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp4 net5 IN4 net3 VDD p12 l = 0.1u w = 0.4u m = 1
mmp5 net5 IN5 VDD VDD p12 l = 0.1u w = 0.21u m = 1


.ends OAI221X2



.subckt OAI222X1 IN1 IN2 IN3 IN4 IN5 IN6 QN VDD VSS
mmp5 net5 IN5 VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp4 net6 IN4 net3 VDD p12 l = 0.1u w = 0.3u m = 1
mmp2 net6 IN2 net1 VDD p12 l = 0.1u w = 0.3u m = 1
mmp6 net6 IN6 net5 VDD p12 l = 0.1u w = 0.3u m = 1
mmp7 net7 net6 VDD VDD p12 l = 0.1u w = 0.37u m = 1
mmp8 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmn5 net6 IN5 net4 VSS n12 l = 0.1u w = 0.14u m = 1
mmn4 net4 IN4 net2 VSS n12 l = 0.1u w = 0.14u m = 1
mmn6 net6 IN6 net4 VSS n12 l = 0.1u w = 0.14u m = 1
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn3 net4 IN3 net2 VSS n12 l = 0.1u w = 0.14u m = 1
mmn7 net7 net6 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn8 QN net7 VSS VSS n12 l = 0.1u w = 0.43u m = 1


.ends OAI222X1



.subckt OAI222X2 IN1 IN2 IN3 IN4 IN5 IN6 QN VDD VSS
mmn5 net6 IN5 net4 VSS n12 l = 0.1u w = 0.14u m = 1
mmn8 QN net7 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmn3 net4 IN3 net2 VSS n12 l = 0.1u w = 0.14u m = 1
mmn4 net4 IN4 net2 VSS n12 l = 0.1u w = 0.14u m = 1
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn7 net7 net6 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn6 net6 IN6 net4 VSS n12 l = 0.1u w = 0.14u m = 1
mmp5 net5 IN5 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp4 net6 IN4 net3 VDD p12 l = 0.1u w = 0.3u m = 1
mmp7 net7 net6 VDD VDD p12 l = 0.1u w = 0.37u m = 1
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp2 net6 IN2 net1 VDD p12 l = 0.1u w = 0.3u m = 1
mmp6 net6 IN6 net5 VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp8 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 2


.ends OAI222X2



.subckt OAI22X1 IN1 IN2 IN3 IN4 QN VDD VSS
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp5 net5 net4 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp4 net4 IN4 net3 VDD p12 l = 0.1u w = 0.5u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp2 net4 IN2 net1 VDD p12 l = 0.1u w = 0.5u m = 1
mmp6 QN net5 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmn3 net4 IN3 net2 VSS n12 l = 0.1u w = 0.23u m = 1
mmn5 net5 net4 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn4 net4 IN4 net2 VSS n12 l = 0.1u w = 0.23u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn6 QN net5 VSS VSS n12 l = 0.1u w = 0.43u m = 1


.ends OAI22X1



.subckt OAI22X2 IN1 IN2 IN3 IN4 QN VDD VSS
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn1 net2 IN1 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn5 net5 net4 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn4 net4 IN4 net2 VSS n12 l = 0.1u w = 0.23u m = 1
mmn3 net4 IN3 net2 VSS n12 l = 0.1u w = 0.23u m = 1
mmn6 QN net5 VSS VSS n12 l = 0.1u w = 0.43u m = 2
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp5 net5 net4 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp6 QN net5 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp4 net4 IN4 net3 VDD p12 l = 0.1u w = 0.5u m = 1
mmp2 net4 IN2 net1 VDD p12 l = 0.1u w = 0.5u m = 1


.ends OAI22X2



.subckt OR2X1 IN1 IN2 Q VDD VSS
mmn2 net1 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 Q net1 VSS VSS n12 l = 0.1u w = 0.48u m = 1
mmn1 net1 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp5 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp2 net2 IN2 VDD VDD p12 l = 0.1u w = 0.9u m = 1
mmp1 net1 IN1 net2 VDD p12 l = 0.1u w = 0.9u m = 1


.ends OR2X1



.subckt OR2X2 IN1 IN2 Q VDD VSS
mmn3 net1 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net1 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 Q net1 VSS VSS n12 l = 0.1u w = 0.48u m = 2
mmp3 net1 IN1 net2 VDD p12 l = 0.1u w = 0.95u m = 1
mmp4 net2 IN2 VDD VDD p12 l = 0.1u w = 0.95u m = 1
mmp6 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 2


.ends OR2X2



.subckt OR2X4 IN1 IN2 Q VDD VSS
mmn3 net1 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net1 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 Q net1 VSS VSS n12 l = 0.1u w = 0.5u m = 4
mmp3 net1 IN1 net2 VDD p12 l = 0.1u w = 0.9u m = 1
mmp4 net2 IN2 VDD VDD p12 l = 0.1u w = 0.9u m = 1
mmp6 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 4


.ends OR2X4



.subckt OR3X1 IN1 IN2 IN3 Q VDD VSS
mmp2 net2 IN2 net3 VDD p12 l = 0.1u w = 1.1u m = 1
mmp5 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp3 net3 IN3 VDD VDD p12 l = 0.1u w = 1.1u m = 1
mmp1 net1 IN1 net2 VDD p12 l = 0.1u w = 1.1u m = 1
mmn1 net1 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net1 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net1 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 Q net1 VSS VSS n12 l = 0.1u w = 0.56u m = 1


.ends OR3X1



.subckt OR3X2 IN1 IN2 IN3 Q VDD VSS
mmn4 net1 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net1 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 Q net1 VSS VSS n12 l = 0.1u w = 0.56u m = 2
mmp6 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp4 net3 IN3 VDD VDD p12 l = 0.1u w = 1.1u m = 1
mmp7 net1 IN1 net2 VDD p12 l = 0.1u w = 1.1u m = 1
mmp8 net2 IN2 net3 VDD p12 l = 0.1u w = 1.1u m = 1


.ends OR3X2



.subckt OR3X4 IN1 IN2 IN3 Q VDD VSS
mmn4 net1 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net1 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 Q net1 VSS VSS n12 l = 0.1u w = 0.64u m = 4
mmp6 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmp4 net3 IN3 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp7 net1 IN1 net2 VDD p12 l = 0.1u w = 1.12u m = 1
mmp8 net2 IN2 net3 VDD p12 l = 0.1u w = 1.12u m = 1


.ends OR3X4



.subckt OR4X1 IN1 IN2 IN3 IN4 Q VDD VSS
mmn5 Q net1 VSS VSS n12 l = 0.1u w = 0.64u m = 1
mmn1 net1 IN1 VSS VSS n12 l = 0.1u w = 0.18u m = 1
mmn4 net1 IN4 VSS VSS n12 l = 0.1u w = 0.18u m = 1
mmn2 net1 IN2 VSS VSS n12 l = 0.1u w = 0.18u m = 1
mmn3 net1 IN3 VSS VSS n12 l = 0.1u w = 0.18u m = 1
mmp1 net1 IN1 net2 VDD p12 l = 0.1u w = 1.12u m = 1
mmp4 net4 IN4 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp5 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp2 net2 IN2 net3 VDD p12 l = 0.1u w = 1.12u m = 1
mmp3 net3 IN3 net4 VDD p12 l = 0.1u w = 1.12u m = 1


.ends OR4X1



.subckt OR4X2 IN1 IN2 IN3 IN4 Q VDD VSS
mmn6 Q net1 VSS VSS n12 l = 0.1u w = 0.64u m = 2
mmn7 net1 IN2 VSS VSS n12 l = 0.1u w = 0.18u m = 1
mmn8 net1 IN1 VSS VSS n12 l = 0.1u w = 0.18u m = 1
mmn9 net1 IN4 VSS VSS n12 l = 0.1u w = 0.18u m = 1
mmn10 net1 IN3 VSS VSS n12 l = 0.1u w = 0.18u m = 1
mmp6 net1 IN1 net2 VDD p12 l = 0.1u w = 1.12u m = 1
mmp7 net4 IN4 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp8 net2 IN2 net3 VDD p12 l = 0.1u w = 1.12u m = 1
mmp9 net3 IN3 net4 VDD p12 l = 0.1u w = 1.12u m = 1
mmp10 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 2


.ends OR4X2



.subckt OR4X4 IN1 IN2 IN3 IN4 Q VDD VSS
mmp6 net1 IN1 net2 VDD p12 l = 0.1u w = 1.12u m = 1
mmp7 net4 IN4 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp8 net2 IN2 net3 VDD p12 l = 0.1u w = 1.12u m = 1
mmp9 net3 IN3 net4 VDD p12 l = 0.1u w = 1.12u m = 1
mmp10 Q net1 VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmn6 Q net1 VSS VSS n12 l = 0.1u w = 0.64u m = 4
mmn7 net1 IN2 VSS VSS n12 l = 0.1u w = 0.16u m = 1
mmn8 net1 IN1 VSS VSS n12 l = 0.1u w = 0.16u m = 1
mmn9 net1 IN4 VSS VSS n12 l = 0.1u w = 0.16u m = 1
mmn10 net1 IN3 VSS VSS n12 l = 0.1u w = 0.16u m = 1


.ends OR4X4



.subckt PGX1 INN INP INQ1 INQ2 VDD VSS
mmp1 INQ1 INP INQ2 VDD p12 l = 0.1u w = 1.12u m = 1
mmn1 INQ1 INN INQ2 VSS n12 l = 0.1u w = 0.35u m = 1


.ends PGX1



.subckt PGX2 INN INP INQ1 INQ2 VDD VSS
mmn1 INQ1 INN INQ2 VSS n12 l = 0.1u w = 0.35u m = 2
mmp1 INQ1 INP INQ2 VDD p12 l = 0.1u w = 1.12u m = 2


.ends PGX2



.subckt PGX4 INN INP INQ1 INQ2 VDD VSS
mmn1 INQ1 INN INQ2 VSS n12 l = 0.1u w = 0.35u m = 4
mmp1 INQ1 INP INQ2 VDD p12 l = 0.1u w = 1.12u m = 4


.ends PGX4



.subckt PMT1 D G S VDD VSS


mg_pmos4t1 D G S VDD p12 l = 0.1u w = 1.12u m = 1
.ends PMT1



.subckt PMT2 D G S VDD VSS
mg_pmos4t1 D G S VDD p12 l = 0.1u w = 1.12u m = 2


.ends PMT2



.subckt PMT3 D G S VDD VSS


mg_pmos4t1 D G S VDD p12 l = 0.1u w = 1.12u m = 4
.ends PMT3



.subckt RDFFARX1 CLK D Q QN RETN RSTB VDD VDDG VSS
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 netp1 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 netp2 D netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 r netp3 VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 netp3 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp7 VDD p12 l = 0.1u w = 0.4u m = 1
mmp7 netp7 CLKN VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp25 netp25 r VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 netp26 netp22 netp25 VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 netp27 netp26 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKP netp27 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 netp5 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp021 r RSTB VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 D netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn7 VSS n12 l = 0.1u w = 0.23u m = 1
mmn8 netn7 CLKP VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.45u m = 1
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 netp26 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 netp26 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp27 netp26 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKN netp27 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn5 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn022 r RSTB VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.22u m = 1


mmp102 netp102 RETNN DL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp101 RETNN RETN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp103 netp103 netp102 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp105 netp102 RETN QL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmn102 netp102 RETN DL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn103 netp103 netp102 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn104 QL netp103 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn105 netp102 RETNN QL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
.ends RDFFARX1



.subckt RDFFARX2 CLK D Q QN RETN RSTB VDD VDDG VSS
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 netp1 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 netp2 D netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 r netp3 VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 netp3 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp7 VDD p12 l = 0.1u w = 0.42u m = 1
mmp7 netp7 CLKN VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp25 netp25 r VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 netp26 netp22 netp25 VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 netp27 netp26 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKP netp27 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 netp5 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp021 r RSTB VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.46u m = 2
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 D netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn7 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 netn7 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 netp26 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 netp26 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp27 netp26 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKN netp27 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn5 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn022 r RSTB VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.22u m = 1


mmp102 netp102 RETNN DL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp101 RETNN RETN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp103 netp103 netp102 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp105 netp102 RETN QL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmn102 netp102 RETN DL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn103 netp103 netp102 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn104 QL netp103 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn105 netp102 RETNN QL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
.ends RDFFARX2



.subckt RDFFNARX1 CLK D Q QN RETN RSTB VDD VDDG VSS


mmn3 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn022 r RSTB VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn8 netn7 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn5 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn7 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 netp26 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 netp26 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp27 netp26 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKP netp27 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 D netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.44u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp2 netp2 D netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp7 VDD p12 l = 0.1u w = 0.55u m = 1
mmp1 netp1 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp5 netp5 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 netp26 netp22 netp25 VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKN netp27 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp3 netp3 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 r netp3 VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 netp7 CLKP VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp27 netp27 netp26 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp021 r RSTB VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp25 netp25 r VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp105 netp102 RETN QL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp101 RETNN RETN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp103 netp103 netp102 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp102 netp102 RETNN DL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmn104 QL netp103 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn102 netp102 RETN DL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn105 netp102 RETNN QL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn103 netp103 netp102 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
.ends RDFFNARX1



.subckt RDFFNARX2 CLK D Q QN RETN RSTB VDD VDDG VSS


mmn3 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn022 r RSTB VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn8 netn7 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn5 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn7 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 netp26 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 netp26 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp27 netp26 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKP netp27 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 D netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.44u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.55u m = 2
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp2 netp2 D netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp7 VDD p12 l = 0.1u w = 0.6u m = 1
mmp1 netp1 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp5 netp5 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 netp26 netp22 netp25 VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKN netp27 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp3 netp3 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 r netp3 VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 netp7 CLKP VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp27 netp27 netp26 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp021 r RSTB VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp25 netp25 r VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp105 netp102 RETN QL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp101 RETNN RETN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp103 netp103 netp102 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp102 netp102 RETNN DL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmn104 QL netp103 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn102 netp102 RETN DL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn105 netp102 RETNN QL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn103 netp103 netp102 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
.ends RDFFNARX2



.subckt RDFFNSRARX1 CLK D NRESTORE Q QN RSTB SAVE VDD VDDG VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 1.1u m = 1
mmp12 net155 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.5u m = 1
mmp7 net155 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net155 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.45u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFNSRARX1



.subckt RDFFNSRARX2 CLK D NRESTORE Q QN RSTB SAVE VDD VDDG VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 1.1u m = 2
mmp12 net155 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.5u m = 2
mmp7 net155 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net155 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.45u m = 2
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.9u m = 2
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFNSRARX2



.subckt RDFFNSRASRNX1 CLK D NRESTORE QN RSTB SAVE SETB VDD VDDG VSS
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net8 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 n20 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp5 net155 RSTB n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 n20 SETB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 n20 _n1 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp16 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net8 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net155 net8 n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 n23 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 _n1 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 _n1 n20 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp14 QN n20 VDD VDD p12 l = 0.1u w = 1.2u m = 1
mmn12 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 n22 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn14 QN n20 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn5 n24 RSTB n25 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 n20 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 n20 _n1 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net5 SETB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net8 n24 VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net8 SETB n22 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net155 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 n25 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 n20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net8 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 _n1 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 _n1 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 _n1 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFNSRASRNX1



.subckt RDFFNSRASRNX2 CLK D NRESTORE QN RSTB SAVE SETB VDD VDDG VSS
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net8 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 n20 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp5 net155 RSTB n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 n20 SETB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 n20 n21 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp16 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net8 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net155 net8 n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 n23 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 n21 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 n21 n20 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp14 QN n20 VDD VDD p12 l = 0.1u w = 1.2u m = 2
mmn12 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 n22 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn14 QN n20 VSS VSS n12 l = 0.1u w = 0.9u m = 2
mmn5 n24 RSTB n25 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 n20 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 n20 n21 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net5 SETB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net8 n24 VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net8 SETB n22 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net155 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 n25 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 n20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net8 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 n21 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 n21 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 n21 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFNSRASRNX2



.subckt RDFFNSRASRQX1 CLK D NRESTORE Q RSTB SAVE SETB VDD VDDG VSS
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net8 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q n21 VDD VDD p12 l = 0.1u w = 1.74u m = 1
mmp12 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 n20 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp5 net155 RSTB n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 n20 SETB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 n20 n21 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp16 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net8 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net155 net8 n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 n23 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 n21 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 n21 n20 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmn12 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 n22 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q n21 VSS VSS n12 l = 0.1u w = 0.69u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn5 n24 RSTB n25 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 n20 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 n20 n21 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net5 SETB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net8 n24 VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net8 SETB n22 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net155 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 n25 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 n20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net8 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 n21 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 n21 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 n21 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFNSRASRQX1



.subckt RDFFNSRASRQX2 CLK D NRESTORE Q RSTB SAVE SETB VDD VDDG VSS
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net8 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q n21 VDD VDD p12 l = 0.1u w = 1.4u m = 2
mmp12 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 n20 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp5 net155 RSTB n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 n20 SETB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 n20 n21 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp16 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net8 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net155 net8 n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 n23 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 n21 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 n21 n20 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmn12 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 n22 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q n21 VSS VSS n12 l = 0.1u w = 0.45u m = 2
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn5 n24 RSTB n25 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 n20 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 n20 n21 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net5 SETB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net8 n24 VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net8 SETB n22 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net155 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 n25 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 n20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net8 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 n21 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 n21 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 n21 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFNSRASRQX2



.subckt RDFFNSRASRX1 CLK D NRESTORE Q QN RSTB SAVE SETB VDD VDDG VSS
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net8 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q n21 VDD VDD p12 l = 0.1u w = 1.3u m = 1
mmp12 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 n20 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp5 net155 RSTB n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 n20 SETB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 n20 n21 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp16 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net8 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net155 net8 n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 n23 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 n21 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 n21 n20 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp14 QN n20 VDD VDD p12 l = 0.1u w = 1.1u m = 1
mmn12 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 n22 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q n21 VSS VSS n12 l = 0.1u w = 0.45u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn14 QN n20 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn5 n24 RSTB n25 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 n20 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 n20 n21 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net5 SETB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net8 n24 VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net8 SETB n22 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net155 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 n25 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 n20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net8 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 n21 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 n21 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 n21 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFNSRASRX1



.subckt RDFFNSRASRX2 CLK D NRESTORE Q QN RSTB SAVE SETB VDD VDDG VSS
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net8 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q n21 VDD VDD p12 l = 0.1u w = 1.25u m = 2
mmp12 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 n20 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp5 net155 RSTB n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 n20 SETB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 n20 n21 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp16 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net8 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net155 net8 n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 n23 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 n21 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 n21 n20 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp14 QN n20 VDD VDD p12 l = 0.1u w = 1.1u m = 2
mmn12 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 n22 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q n21 VSS VSS n12 l = 0.1u w = 0.45u m = 2
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn14 QN n20 VSS VSS n12 l = 0.1u w = 0.9u m = 2
mmn5 n24 RSTB n25 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 n20 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 n20 n21 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net5 SETB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net8 n24 VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net8 SETB n22 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net155 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 n25 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 n20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net8 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 n21 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 n21 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 n21 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFNSRASRX2



.subckt RDFFNSRASX1 CLK D NRESTORE Q QN SAVE SETB VDD VDDG VSS
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net8 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q n21 VDD VDD p12 l = 0.1u w = 1.3u m = 1
mmp12 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 n20 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp5 net155 VDD n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 n20 SETB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 n20 n21 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp16 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net8 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net155 net8 n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 n23 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 n21 VDD VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 n21 n20 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp14 QN n20 VDD VDD p12 l = 0.1u w = 1.1u m = 1
mmn12 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 n22 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q n21 VSS VSS n12 l = 0.1u w = 0.45u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn14 QN n20 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn5 n24 VDD n25 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 n20 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 n20 n21 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net5 SETB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net8 n24 VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net8 SETB n22 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net155 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 n25 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 n20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net8 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 n21 VDD net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 n21 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 n21 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFNSRASX1



.subckt RDFFNSRASX2 CLK D NRESTORE Q QN SAVE SETB VDD VDDG VSS
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net8 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q n21 VDD VDD p12 l = 0.1u w = 1.25u m = 2
mmp12 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 n20 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp5 net155 VDD n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 n20 SETB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 n20 n21 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp16 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net8 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net155 net8 n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 n23 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 n21 VDD VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 n21 n20 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp14 QN n20 VDD VDD p12 l = 0.1u w = 1.1u m = 2
mmn12 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 n22 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q n21 VSS VSS n12 l = 0.1u w = 0.45u m = 2
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn14 QN n20 VSS VSS n12 l = 0.1u w = 0.9u m = 2
mmn5 n24 VDD n25 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 n20 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 n20 n21 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net5 SETB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net8 n24 VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net8 SETB n22 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net155 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 n25 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 n20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net8 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 n21 VDD net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 n21 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 n21 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFNSRASX2



.subckt RDFFNSRX1 CLK D NRESTORE Q QN SAVE VDD VDDG VSS
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 1u m = 1
mmp12 net155 net8 net1000 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp60 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net1000 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKN hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.6u m = 1
mmp7 net155 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp61 net1 net2 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp03 hjf D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn1 net1 CLKP hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn60 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn61 net1 net2 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net155 net8 net1222 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.6u m = 1
mmn8 net8 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.6u m = 1
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net1222 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn03 hjf D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1


.ends RDFFNSRX1



.subckt RDFFNSRX2 CLK D NRESTORE Q QN SAVE VDD VDDG VSS
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 0.8u m = 2
mmp12 net155 net8 net1000 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp60 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net1000 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKN hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.64u m = 2
mmp7 net155 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp61 net1 net2 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp03 hjf D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn1 net1 CLKP hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn60 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn61 net1 net2 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net155 net8 net1222 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.6u m = 2
mmn8 net8 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.59u m = 2
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net1222 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn03 hjf D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1


.ends RDFFNSRX2



.subckt RDFFNX1 CLK D Q QN RETN VDD VDDG VSS
mmp26 netp25 netp22 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 netp1 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 netp2 D netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp6 VDD p12 l = 0.1u w = 0.56u m = 1
mmp7 netp6 CLKP VDD VDD p12 l = 0.1u w = 0.56u m = 1
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp27 netp26 netp25 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKN netp26 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 netp5 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp103 netp103 netp102 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp105 netp102 RETN QL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp102 netp102 RETNN DL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp101 RETNN RETN VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmn26 netp25 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 D netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 netn6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp26 netp25 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKP netp26 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn4 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.44u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn103 netp103 netp102 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn104 QL netp103 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn105 netp102 RETNN QL VSS n12 l = 0.1u w = 0.21u m = 1
mmn102 netp102 RETN DL VSS n12 l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends RDFFNX1



.subckt RDFFNX2 CLK D Q QN RETN VDD VDDG VSS
mmp26 netp25 netp22 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 netp1 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 netp2 D netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp6 VDD p12 l = 0.1u w = 0.65u m = 1
mmp7 netp6 CLKP VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp27 netp26 netp25 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKN netp26 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 netp5 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp103 netp103 netp102 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp105 netp102 RETN QL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp102 netp102 RETNN DL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp101 RETNN RETN VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmn26 netp25 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.55u m = 2
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 D netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn6 VSS n12 l = 0.1u w = 0.23u m = 1
mmn8 netn6 CLKN VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp26 netp25 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKP netp26 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn4 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn103 netp103 netp102 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn104 QL netp103 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn105 netp102 RETNN QL VSS n12 l = 0.1u w = 0.21u m = 1
mmn102 netp102 RETN DL VSS n12 l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends RDFFNX2



.subckt RDFFSRARX1 CLK D NRESTORE Q QN RSTB SAVE VDD VDDG VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net2 RESTORE aa VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp19 aa jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net155 CLKN aa VDD p12 l = 0.1u w = 0.45u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 1.1u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.5u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net155 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net2 NRESTORE aa VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn18 aa jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKP aa VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn12 net155 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.45u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFSRARX1



.subckt RDFFSRARX2 CLK D NRESTORE Q QN RSTB SAVE VDD VDDG VSS
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net2 RESTORE aa VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp19 aa jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net155 CLKN aa VDD p12 l = 0.1u w = 0.45u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 0.9u m = 2
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.5u m = 2
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net155 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net2 NRESTORE aa VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn18 aa jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKP aa VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.9u m = 2
mmn12 net155 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.35u m = 2
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFSRARX2



.subckt RDFFSRASRX1 CLK D NRESTORE Q QN RSTB SAVE SETB VDD VDDG VSS
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net8 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q n21 VDD VDD p12 l = 0.1u w = 1.3u m = 1
mmp12 net2564 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 n20 CLKN _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp5 net155 RSTB n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 n20 SETB net2564 VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 n20 n21 net2564 VDD p12 l = 0.1u w = 0.33u m = 1
mmp16 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net8 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net155 net8 n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 n23 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 n21 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 n21 n20 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp14 QN n20 VDD VDD p12 l = 0.1u w = 1.1u m = 1
mmn12 _n11 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 n22 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q n21 VSS VSS n12 l = 0.1u w = 0.45u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn14 QN n20 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn5 n24 RSTB n25 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 n20 CLKP _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 n20 n21 _n8 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n8 SETB _n11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net8 n24 VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net8 SETB n22 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net155 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 n25 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 n20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net8 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 n21 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 n21 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 n21 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFSRASRX1



.subckt RDFFSRASRX2 CLK D NRESTORE Q QN RSTB SAVE SETB VDD VDDG VSS
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net8 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q n21 VDD VDD p12 l = 0.1u w = 1.3u m = 2
mmp12 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 n20 CLKN _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp5 net155 RSTB n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 n20 SETB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 n20 n21 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp16 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net8 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net155 net8 n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 n23 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 n21 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 n21 n20 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp14 QN n20 VDD VDD p12 l = 0.1u w = 1.1u m = 2
mmn12 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 n22 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q n21 VSS VSS n12 l = 0.1u w = 0.45u m = 2
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn14 QN n20 VSS VSS n12 l = 0.1u w = 0.9u m = 2
mmn5 n24 RSTB n25 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 n20 CLKP _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 n20 n21 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net5 SETB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net8 n24 VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net8 SETB n22 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net155 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 n25 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 n20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net8 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 n21 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 n21 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 n21 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFSRASRX2



.subckt RDFFSRASX1 CLK D NRESTORE Q QN SAVE SETB VDD VDDG VSS
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net8 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q n21 VDD VDD p12 l = 0.1u w = 1.3u m = 1
mmp12 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 n20 CLKN _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp5 net155 VDD n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 n20 SETB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 n20 n21 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp16 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net8 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net155 net8 n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 n23 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 n21 VDD VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 n21 n20 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp14 QN n20 VDD VDD p12 l = 0.1u w = 1.1u m = 1
mmn12 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 n22 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q n21 VSS VSS n12 l = 0.1u w = 0.45u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn14 QN n20 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn5 n24 VDD n25 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 n20 CLKP _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 n20 n21 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net5 SETB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net8 n24 VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net8 SETB n22 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net155 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 n25 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 n20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net8 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 n21 VDD net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 n21 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 n21 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFSRASX1



.subckt RDFFSRASX2 CLK D NRESTORE Q QN SAVE SETB VDD VDDG VSS
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net8 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp13 Q n21 VDD VDD p12 l = 0.1u w = 1.3u m = 2
mmp12 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 n20 CLKN _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp5 net155 VDD n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 n20 SETB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 n20 n21 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp16 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp03 net06 D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net8 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net155 net8 n23 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 n23 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 n21 VDD VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp8 n21 n20 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp14 QN n20 VDD VDD p12 l = 0.1u w = 1.1u m = 2
mmn12 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 n22 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q n21 VSS VSS n12 l = 0.1u w = 0.45u m = 2
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn14 QN n20 VSS VSS n12 l = 0.1u w = 0.9u m = 2
mmn5 n24 VDD n25 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 n20 CLKP _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 n20 n21 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net5 SETB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net8 n24 VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net8 SETB n22 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net155 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 n25 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 n20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net8 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 n21 VDD net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 n21 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 n21 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFSRASX2



.subckt RDFFSRSSRX1 CLK D NRESTORE Q QN RSTB SAVE SETB VDD VDDG VSS
mmp03 net06 net0666 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net2 RESTORE aa VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp19 aa jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net155 CLKN aa VDD p12 l = 0.1u w = 0.45u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp14 Q net155 VDD VDD p12 l = 0.1u w = 1.1u m = 1
mmp13 QN net8 VDD VDD p12 l = 0.1u w = 1.5u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 VDD VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp5 net1 VDD net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net155 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 SET SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp16 net0666 D net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net0666 RSTB net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 net01 SET VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn03 net06 net0666 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net2 NRESTORE aa VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 VDD net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn18 aa jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKP aa VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 Q net155 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn12 net155 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 VDD net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 QN net8 VSS VSS n12 l = 0.1u w = 0.45u m = 1
mmn3 SET SETB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net03 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 net0666 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net0666 SET net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFSRSSRX1



.subckt RDFFSRSSRX2 CLK D NRESTORE Q QN RSTB SAVE SETB VDD VDDG VSS
mmp03 net06 net0678 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net2 RESTORE aa VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp19 aa jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net155 CLKN aa VDD p12 l = 0.1u w = 0.45u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp14 Q net155 VDD VDD p12 l = 0.1u w = 0.9u m = 2
mmp13 QN net8 VDD VDD p12 l = 0.1u w = 1.5u m = 2
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 VDD VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp5 net1 VDD net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net155 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 SET SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp16 net0678 RSTB net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net0678 D net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 net01 SET VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn03 net06 net0678 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net2 NRESTORE aa VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 VDD net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn18 aa jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKP aa VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 Q net155 VSS VSS n12 l = 0.1u w = 0.9u m = 2
mmn12 net155 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 VDD net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 QN net8 VSS VSS n12 l = 0.1u w = 0.35u m = 2
mmn3 SET SETB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net0678 SET net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 net0678 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net03 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RDFFSRSSRX2



.subckt RDFFSRX1 CLK D NRESTORE Q QN SAVE VDD VDDG VSS
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 1u m = 1
mmp12 net155 net8 net1000 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp60 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net1000 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.6u m = 1
mmp7 net155 CLKN _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp61 net1 net2 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp03 hjf D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn1 net1 CLKN hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKP _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn60 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn61 net1 net2 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net155 net8 net1222 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.6u m = 1
mmn8 net8 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.6u m = 1
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net1222 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn03 hjf D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1


.ends RDFFSRX1



.subckt RDFFSRX2 CLK D NRESTORE Q QN SAVE VDD VDDG VSS
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 0.8u m = 2
mmp12 net155 net8 net1000 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp60 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net1000 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.64u m = 2
mmp7 net155 CLKN _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp61 net1 net2 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp03 hjf D VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn1 net1 CLKN hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKP _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn60 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn61 net1 net2 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net155 net8 net1222 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.6u m = 2
mmn8 net8 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.59u m = 2
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net1222 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn03 hjf D VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1


.ends RDFFSRX2



.subckt RDFFX1 CLK D Q QN RETN VDD VDDG VSS
mmp26 netp25 netp22 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 netp1 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 netp2 D netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp6 VDD p12 l = 0.1u w = 0.41u m = 1
mmp7 netp6 CLKN VDD VDD p12 l = 0.1u w = 0.41u m = 1
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp27 netp26 netp25 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKP netp26 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 netp5 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp103 netp103 netp102 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp105 netp102 RETN QL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp102 netp102 RETNN DL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp101 RETNN RETN VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmn26 netp25 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 D netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn6 VSS n12 l = 0.1u w = 0.23u m = 1
mmn8 netn6 CLKP VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp26 netp25 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKN netp26 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn4 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn103 netp103 netp102 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn104 QL netp103 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn105 netp102 RETNN QL VSS n12 l = 0.1u w = 0.21u m = 1
mmn102 netp102 RETN DL VSS n12 l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends RDFFX1



.subckt RDFFX2 CLK D Q QN RETN VDD VDDG VSS
mmp26 netp25 netp22 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 netp1 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 netp2 D netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp6 VDD p12 l = 0.1u w = 0.45u m = 1
mmp7 netp6 CLKN VDD VDD p12 l = 0.1u w = 0.45u m = 1
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp27 netp26 netp25 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKP netp26 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 netp5 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp103 netp103 netp102 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp105 netp102 RETN QL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp102 netp102 RETNN DL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp101 RETNN RETN VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmn26 netp25 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.46u m = 2
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 D netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 netn6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp26 netp25 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKN netp26 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn4 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn103 netp103 netp102 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn104 QL netp103 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn105 netp102 RETNN QL VSS n12 l = 0.1u w = 0.21u m = 1
mmn102 netp102 RETN DL VSS n12 l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends RDFFX2



.subckt RSDFFARX1 CLK D Q QN RETN RSTB SE SI VDD VDDG VSS
mmp03 INN D netp02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 netp04 netp01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 INN SI netp04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp01 netp01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 netp02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 netp1 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 netp2 INP netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 r netp3 VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 netp3 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp7 VDD p12 l = 0.1u w = 0.37u m = 1
mmp7 netp7 CLKN VDD VDD p12 l = 0.1u w = 0.37u m = 1
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp25 netp25 r VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 netp26 netp22 netp25 VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 netp27 netp26 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKP netp27 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 netp5 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp021 r RSTB VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp06 INP INN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 netp01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 INN SI netn04 VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 netn04 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 netn02 netp01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 INN D netn02 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 INP netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn7 VSS n12 l = 0.1u w = 0.23u m = 1
mmn8 netn7 CLKP VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.45u m = 1
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 netp26 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 netp26 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp27 netp26 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKN netp27 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn5 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn022 r RSTB VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn06 INP INN VSS VSS n12 l = 0.1u w = 0.21u m = 1



mmp101 RETNN RETN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp103 netp103 netp102 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp105 netp102 RETN QL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp102 netp102 RETNN DL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmn102 netp102 RETN DL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn103 netp103 netp102 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn104 QL netp103 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn105 netp102 RETNN QL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
.ends RSDFFARX1



.subckt RSDFFARX2 CLK D Q QN RETN RSTB SE SI VDD VDDG VSS
mmp03 INN D netp02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 netp04 netp01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 INN SI netp04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp01 netp01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 netp02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 netp1 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 netp2 INP netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 r netp3 VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 netp3 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp7 VDD p12 l = 0.1u w = 0.44u m = 1
mmp7 netp7 CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp25 netp25 r VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 netp26 netp22 netp25 VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 netp27 netp26 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKP netp27 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 netp5 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp021 r RSTB VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp06 INP INN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 netp01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 INN SI netn04 VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 netn04 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 netn02 netp01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 INN D netn02 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.44u m = 2
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 INP netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn7 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 netn7 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 netp26 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 netp26 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp27 netp26 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKN netp27 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn5 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn022 r RSTB VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn06 INP INN VSS VSS n12 l = 0.1u w = 0.21u m = 1



mmp105 netp102 RETN QL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp102 netp102 RETNN DL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp101 RETNN RETN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp103 netp103 netp102 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmn105 netp102 RETNN QL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn102 netp102 RETN DL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn103 netp103 netp102 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn104 QL netp103 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
.ends RSDFFARX2



.subckt RSDFFNARX1 CLK D Q QN RETN RSTB SE SI VDD VDDG VSS
mmp03 INN D netp02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 netp04 netp01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 INN SI netp04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp01 netp01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 netp02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 netp1 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 netp2 INP netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 r netp3 VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 netp3 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp7 VDD p12 l = 0.1u w = 0.55u m = 1
mmp7 netp7 CLKP VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp25 netp25 r VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 netp26 netp22 netp25 VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 netp27 netp26 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKN netp27 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 netp5 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp021 r RSTB VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp06 INP INN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 netp01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 INN SI netn04 VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 netn04 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 netn02 netp01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 INN D netn02 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.55u m = 1
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 INP netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn7 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 netn7 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 netp26 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 netp26 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp27 netp26 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKP netp27 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn5 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn022 r RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.44u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn06 INP INN VSS VSS n12 l = 0.1u w = 0.21u m = 1



mmp101 RETNN RETN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp103 netp103 netp102 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp105 netp102 RETN QL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp102 netp102 RETNN DL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmn102 netp102 RETN DL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn103 netp103 netp102 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn104 QL netp103 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn105 netp102 RETNN QL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
.ends RSDFFNARX1



.subckt RSDFFNARX2 CLK D Q QN RETN RSTB SE SI VDD VDDG VSS
mmp03 INN D netp02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 netp04 netp01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 INN SI netp04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp01 netp01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 netp02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 netp1 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 netp2 INP netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 r netp3 VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 netp3 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp7 VDD p12 l = 0.1u w = 0.6u m = 1
mmp7 netp7 CLKP VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp25 netp25 r VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 netp26 netp22 netp25 VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 netp27 netp26 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKN netp27 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 netp5 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp021 r RSTB VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp06 INP INN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 netp01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 INN SI netn04 VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 netn04 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 netn02 netp01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 INN D netn02 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.55u m = 2
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 INP netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn7 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 netn7 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 netp26 r VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 netp26 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp27 netp26 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKP netp27 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn5 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn022 r RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.44u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn06 INP INN VSS VSS n12 l = 0.1u w = 0.21u m = 1



mmp105 netp102 RETN QL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp102 netp102 RETNN DL VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp101 RETNN RETN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp103 netp103 netp102 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmn105 netp102 RETNN QL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn102 netp102 RETN DL VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn103 netp103 netp102 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn104 QL netp103 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
.ends RSDFFNARX2



.subckt RSDFFNSRARX1 CLK D NRESTORE Q QN RSTB SAVE SE SI VDD VDDG VSS
mmp23 rrr _n53 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp12 net155 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKN hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.68u m = 1
mmp7 net155 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp3 _n50 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 _n53 D _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5 p1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 hjf rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 p1 SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 _n53 SI net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmn24 rrr _n53 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net1 CLKP hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 _n991 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 _n989 RSTB _n991 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net155 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.44u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 _n989 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.46u m = 1
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 _n52 p1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 _n53 SI net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n53 D _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 hjf rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 p1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFNSRARX1



.subckt RSDFFNSRARX2 CLK D NRESTORE Q QN RSTB SAVE SE SI VDD VDDG VSS
mmp03 net06 rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 0.58u m = 2
mmp12 net155 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.56u m = 2
mmp7 net155 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp3 net2m SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 net3m D net2m VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5m net1m VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp23 rrr net3m VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp24 net1m SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 net3m SI net5m VDD p12 l = 0.1u w = 0.65u m = 1
mmn03 net06 rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net155 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.44u m = 2
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.41u m = 2
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 net4m net1m VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6m SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 net3m SI net6m VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net3m D net4m VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 rrr net3m VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn25 net1m SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFNSRARX2



.subckt RSDFFNSRASRNX1 CLK D NRESTORE QN RSTB SAVE SE SETB SI VDD VDDG VSS
mmp23 rrr _n53 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp14 QN net1556 VDD VDD p12 l = 0.1u w = 0.9u m = 1
mmp10 net444 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 net2 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net1556 net8 net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net1556 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 net2 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net1556 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net155 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp29 net1556 SETB net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net155 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 _n50 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 _n53 D _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5 p1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 hjf rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 p1 SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 _n53 SI net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmn24 rrr _n53 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net155 CLKP hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net1556 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 _n991 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 net2 SETB net994 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 _n989 RSTB _n991 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 _n1248 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 net994 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net1556 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 _n1247 SETB _n1248 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net2 _n989 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net1556 VSS VSS n12 l = 0.1u w = 0.46u m = 1
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn29 net1556 net8 _n1247 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 _n52 p1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 _n53 SI net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n53 D _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 hjf rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 p1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFNSRASRNX1



.subckt RSDFFNSRASRNX2 CLK D NRESTORE QN RSTB SAVE SE SETB SI VDD VDDG VSS
mmp23 rrr _n53 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp14 QN net1556 VDD VDD p12 l = 0.1u w = 0.96u m = 2
mmp10 net444 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 net2 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net1556 net8 net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net1556 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 net2 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net1556 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net155 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp29 net1556 SETB net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net155 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 _n50 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 _n53 D _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5 p1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 hjf rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 p1 SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 _n53 SI net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmn24 rrr _n53 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net155 CLKP hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net1556 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 _n991 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 net2 SETB net994 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 _n989 RSTB _n991 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 _n1248 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 net994 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net1556 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 _n1247 SETB _n1248 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net2 _n989 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net1556 VSS VSS n12 l = 0.1u w = 0.59u m = 2
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn29 net1556 net8 _n1247 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 _n52 p1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 _n53 SI net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n53 D _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 hjf rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 p1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFNSRASRNX2



.subckt RSDFFNSRASRQX1 CLK D NRESTORE Q RSTB SAVE SE SETB SI VDD VDDG VSS
mmp23 rrr _n53 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp10 net444 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 net2 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net1556 net8 net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.4u m = 1
mmp7 net1556 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 net2 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net1556 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net155 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp29 net1556 SETB net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net155 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 _n50 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 _n53 D _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5 p1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 hjf rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 p1 SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 _n53 SI net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmn24 rrr _n53 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net155 CLKP hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net1556 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 _n991 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 net2 SETB net994 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 _n989 RSTB _n991 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 _n1248 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.81u m = 1
mmn28 net994 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net1556 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 _n1247 SETB _n1248 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net2 _n989 VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn29 net1556 net8 _n1247 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 _n52 p1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 _n53 SI net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n53 D _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 hjf rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 p1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFNSRASRQX1



.subckt RSDFFNSRASRQX2 CLK D NRESTORE Q RSTB SAVE SE SETB SI VDD VDDG VSS
mmp23 rrr _n53 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp10 net444 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 net2 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net1556 net8 net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.1u m = 2
mmp7 net1556 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 net2 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net1556 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net155 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp29 net1556 SETB net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net155 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 _n50 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 _n53 D _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5 p1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 hjf rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 p1 SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 _n53 SI net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmn24 rrr _n53 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net155 CLKP hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net1556 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 _n991 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 net2 SETB net994 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 _n989 RSTB _n991 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 _n1248 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.81u m = 2
mmn28 net994 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net1556 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 _n1247 SETB _n1248 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net2 _n989 VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn29 net1556 net8 _n1247 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 _n52 p1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 _n53 SI net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n53 D _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 hjf rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 p1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFNSRASRQX2



.subckt RSDFFNSRASRX1 CLK D NRESTORE Q QN RSTB SAVE SE SETB SI VDD VDDG VSS
mmp23 rrr _n53 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp14 QN net1556 VDD VDD p12 l = 0.1u w = 0.75u m = 1
mmp10 net444 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 net2 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net1556 net8 net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.7u m = 1
mmp7 net1556 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 net2 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net1556 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net155 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp29 net1556 SETB net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net155 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 _n50 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 _n53 D _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5 p1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 hjf rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 p1 SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 _n53 SI net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmn24 rrr _n53 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net155 CLKP hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net1556 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 _n991 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 net2 SETB net994 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 _n989 RSTB _n991 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 _n1248 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.55u m = 1
mmn28 net994 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net1556 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 _n1247 SETB _n1248 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net2 _n989 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net1556 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn29 net1556 net8 _n1247 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 _n52 p1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 _n53 SI net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n53 D _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 hjf rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 p1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFNSRASRX1



.subckt RSDFFNSRASRX2 CLK D NRESTORE Q QN RSTB SAVE SE SETB SI VDD VDDG VSS
mmp23 rrr _n53 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp14 QN net1556 VDD VDD p12 l = 0.1u w = 0.75u m = 2
mmp10 net444 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 net2 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net1556 net8 net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.7u m = 2
mmp7 net1556 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 net2 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net1556 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net155 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp29 net1556 SETB net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net155 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 _n50 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 _n53 D _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5 p1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 hjf rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 p1 SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 _n53 SI net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmn24 rrr _n53 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net155 CLKP hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net1556 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 _n991 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 net2 SETB net994 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 _n989 RSTB _n991 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 _n1248 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn28 net994 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net1556 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 _n1247 SETB _n1248 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net2 _n989 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net1556 VSS VSS n12 l = 0.1u w = 0.46u m = 2
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn29 net1556 net8 _n1247 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 _n52 p1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 _n53 SI net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n53 D _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 hjf rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 p1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFNSRASRX2



.subckt RSDFFNSRASX1 CLK D NRESTORE Q QN SAVE SE SETB SI VDD VDDG VSS
mmp23 rrr _n53 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp14 QN net1556 VDD VDD p12 l = 0.1u w = 0.75u m = 1
mmp10 net444 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 net2 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net1556 net8 net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.7u m = 1
mmp7 net1556 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 net2 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net1556 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net155 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp29 net1556 SETB net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net155 VDD net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 VDD VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 _n50 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 _n53 D _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5 p1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 hjf rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 p1 SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 _n53 SI net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmn24 rrr _n53 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net155 CLKP hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net1556 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 _n991 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 net2 SETB net994 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 _n989 VDD _n991 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 _n1248 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.55u m = 1
mmn28 net994 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 VDD net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net1556 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 _n1247 SETB _n1248 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net2 _n989 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net1556 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn29 net1556 net8 _n1247 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 _n52 p1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 _n53 SI net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n53 D _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 hjf rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 p1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFNSRASX1



.subckt RSDFFNSRASX2 CLK D NRESTORE Q QN SAVE SE SETB SI VDD VDDG VSS
mmp23 rrr _n53 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp14 QN net1556 VDD VDD p12 l = 0.1u w = 0.75u m = 2
mmp10 net444 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 net2 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net1556 net8 net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKN hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.7u m = 2
mmp7 net1556 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 net2 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net1556 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net155 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp29 net1556 SETB net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net155 VDD net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 VDD VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 _n50 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 _n53 D _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5 p1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 hjf rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 p1 SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 _n53 SI net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmn24 rrr _n53 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net155 CLKP hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net1556 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 _n991 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 net2 SETB net994 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 _n989 VDD _n991 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 _n1248 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn28 net994 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 VDD net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net1556 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 _n1247 SETB _n1248 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net2 _n989 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net1556 VSS VSS n12 l = 0.1u w = 0.46u m = 2
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn29 net1556 net8 _n1247 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 _n52 p1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 _n53 SI net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n53 D _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 hjf rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 p1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFNSRASX2



.subckt RSDFFNSRX1 CLK D NRESTORE Q QN SAVE SE SI VDD VDDG VSS
mmp23 rrr _n53 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 0.8u m = 1
mmp12 net155 net8 net1000 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp60 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net1000 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKN hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.64u m = 1
mmp7 net155 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp61 net1 net2 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 _n50 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 _n53 D _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5 p1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 hjf rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 p1 SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 _n53 SI net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmn24 rrr _n53 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net1 CLKP hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn60 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn61 net1 net2 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net155 net8 net1222 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.6u m = 1
mmn8 net8 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.6u m = 1
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net1222 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 _n52 p1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 _n53 SI net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n53 D _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 hjf rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 p1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFNSRX1



.subckt RSDFFNSRX2 CLK D NRESTORE Q QN SAVE SE SI VDD VDDG VSS
mmp23 rrr _n53 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 0.8u m = 2
mmp12 net155 net8 net1000 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp60 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net1000 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKN hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.6u m = 2
mmp7 net155 CLKP _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp61 net1 net2 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 _n50 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 _n53 D _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5 p1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 hjf rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 p1 SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 _n53 SI net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmn24 rrr _n53 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net1 CLKP hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKN _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn60 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn61 net1 net2 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net155 net8 net1222 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.6u m = 2
mmn8 net8 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.59u m = 2
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net1222 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 _n52 p1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 _n53 SI net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n53 D _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 hjf rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 p1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFNSRX2



.subckt RSDFFNX1 CLK D Q QN RETN SE SI VDD VDDG VSS
mmp26 netp26 netp22 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 netp02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp01 netp01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 INN SI netp04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp06 INP INN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 netp1 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 netp2 INP netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 INN D netp02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp6 VDD p12 l = 0.1u w = 0.57u m = 1
mmp7 netp6 CLKP VDD VDD p12 l = 0.1u w = 0.57u m = 1
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp04 netp04 netp01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 netp27 netp26 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKN netp27 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 netp5 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp103 netp103 netp102 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp105 netp102 RETN QL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp102 netp102 RETNN DL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp101 RETNN RETN VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmn26 netp26 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn06 INP INN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 netn02 netp01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 INN SI netn04 VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 netn04 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 INP netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 INN D netn02 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 netn6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 netp01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp27 netp26 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKP netp27 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn5 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.44u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn103 netp103 netp102 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn104 QL netp103 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn105 netp102 RETNN QL VSS n12 l = 0.1u w = 0.21u m = 1
mmn102 netp102 RETN DL VSS n12 l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends RSDFFNX1



.subckt RSDFFNX2 CLK D Q QN RETN SE SI VDD VDDG VSS
mmp26 netp26 netp22 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 netp02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp01 netp01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 INN SI netp04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp06 INP INN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 netp1 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 netp2 INP netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 INN D netp02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp6 VDD p12 l = 0.1u w = 0.6u m = 1
mmp7 netp6 CLKP VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp04 netp04 netp01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 netp27 netp26 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKN netp27 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 netp5 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp103 netp103 netp102 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp105 netp102 RETN QL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp102 netp102 RETNN DL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp101 RETNN RETN VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmn26 netp26 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn06 INP INN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 netn02 netp01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 INN SI netn04 VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 netn04 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.55u m = 2
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 INP netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 INN D netn02 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 netn6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 netp01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp27 netp26 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKP netp27 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn5 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.44u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn103 netp103 netp102 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn104 QL netp103 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn105 netp102 RETNN QL VSS n12 l = 0.1u w = 0.21u m = 1
mmn102 netp102 RETN DL VSS n12 l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends RSDFFNX2



.subckt RSDFFSRARX1 CLK D NRESTORE Q QN RSTB SAVE SE SI VDD VDDG VSS
mmn15 jk for_t VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 for_t jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 for_t net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk for_t VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 for_t jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 for_t net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp24 _n2 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp23 nn1 D _n2 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 _n50 nn VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 nn1 SI _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp25 ff nn1 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp3 nn SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp03 net06 ff VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net155 CLKN _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp12 net155 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.25u m = 1
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 0.9u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmn25 nn1 D _n4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n4 nn VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 nn1 SI _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 _n52 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 ff nn1 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn3 nn SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net06 ff VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKP _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net155 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
.ends RSDFFSRARX1



.subckt RSDFFSRARX2 CLK D NRESTORE Q QN RSTB SAVE SE SI VDD VDDG VSS
mmp03 net06 ff VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 0.8u m = 2
mmp12 net155 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.5u m = 2
mmp7 net155 CLKN _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 ff nn1 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp16 nn1 SI _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp24 _n2 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp3 nn SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp23 nn1 D _n2 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 _n50 nn VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmn03 net06 ff VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKP _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net155 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.35u m = 2
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.8u m = 2
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn17 ff nn1 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn25 nn1 D _n4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 _n52 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 nn1 SI _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 nn SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n4 nn VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFSRARX2



.subckt RSDFFSRASRX1 CLK D NRESTORE Q QN RSTB SAVE SE SETB SI VDD VDDG VSS
mmp23 rrr _n53 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp14 QN net1556 VDD VDD p12 l = 0.1u w = 1.18u m = 1
mmp10 net444 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 net2 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net1556 net8 net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKP hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.18u m = 1
mmp7 net1556 CLKN _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 net2 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net1556 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net155 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp29 net1556 SETB net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net155 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 _n50 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 _n53 D _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5 p1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 hjf rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 p1 SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 _n53 SI net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmn24 rrr _n53 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net155 CLKN hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net1556 CLKP _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 _n991 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 net2 SETB net994 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 _n989 RSTB _n991 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 _n1248 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.46u m = 1
mmn28 net994 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net1556 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 _n1247 SETB _n1248 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net2 _n989 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net1556 VSS VSS n12 l = 0.1u w = 0.46u m = 1
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn29 net1556 net8 _n1247 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 _n52 p1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 _n53 SI net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n53 D _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 hjf rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 p1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1


.ends RSDFFSRASRX1



.subckt RSDFFSRASRX2 CLK D NRESTORE Q QN RSTB SAVE SE SETB SI VDD VDDG VSS
mmp23 rrr _n53 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp14 QN net1556 VDD VDD p12 l = 0.1u w = 1.18u m = 2
mmp10 net444 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 net2 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net1556 net8 net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net155 CLKP hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.18u m = 2
mmp7 net1556 CLKN _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 net2 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net1556 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp6 net155 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp29 net1556 SETB net444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net155 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 _n50 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 _n53 D _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5 p1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 hjf rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 p1 SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 _n53 SI net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmn24 rrr _n53 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net155 CLKN hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net1556 CLKP _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 _n991 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 net2 SETB net994 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 _n989 RSTB _n991 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 _n1248 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.48u m = 2
mmn28 net994 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net1556 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 _n1247 SETB _n1248 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net155 net2 _n989 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net1556 VSS VSS n12 l = 0.1u w = 0.48u m = 2
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn29 net1556 net8 _n1247 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 _n52 p1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 _n53 SI net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n53 D _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 hjf rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 p1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1


.ends RSDFFSRASRX2



.subckt RSDFFSRASX1 CLK D NRESTORE Q QN SAVE SE SETB SI VDD VDDG VSS
mmn28 aa jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 nn SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.52u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKP aa VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net06 net_146 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net112589 SETB Mushegh VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn29 QN net155 VSS VSS n12 l = 0.1u w = 0.52u m = 1
mmn12 Mushegh net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 nn1 D _n2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 VDD net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 net_146 nn1 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn23 _n2 nn VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 nn1 SI _n3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 _n3 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net112589 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net112589 NRESTORE aa VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 VDD net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn30 net155 net8 net5555555 VSS n12 l = 0.1u w = 0.21u m = 1
mmn31 net5555555 SETB net6666666 VSS n12 l = 0.1u w = 0.21u m = 1
mmn34 net6666666 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp13 net06 net_146 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 net112589 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp12 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp3 nn SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp27 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp25 net_146 nn1 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp6 net1 net112589 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 aa jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 0.8u m = 1
mmp5 net1 VDD net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp23 nn1 D _n1 VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 nn1 SI _n4 VDD p12 l = 0.1u w = 0.65u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp21 Q net8 VDD VDD p12 l = 0.1u w = 1.56u m = 1
mmp7 net155 CLKN aa VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net112589 RESTORE aa VDD p12 l = 0.1u w = 0.33u m = 1
mmp29 net112589 net1 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp24 _n1 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp9 net8 VDD VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp17 _n4 nn VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp30 net444444 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp31 net155 SETB net444444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp34 net155 net8 net444444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp28 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
.ends RSDFFSRASX1



.subckt RSDFFSRASX2 CLK D NRESTORE Q QN SAVE SE SETB SI VDD VDDG VSS
mmn30 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn31 net06 net_146 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn34 net8 VDD net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn35 _n7 nn VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn36 net5 VDD net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn37 net112589 SETB Mushegh VSS n12 l = 0.1u w = 0.21u m = 1
mmn39 net155 CLKP aa VSS n12 l = 0.1u w = 0.21u m = 1
mmn40 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn41 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn42 net_146 nn1 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn44 net6666666 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn45 QN net155 VSS VSS n12 l = 0.1u w = 0.96u m = 1
mmn47 net1 net112589 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn49 net9 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn51 Q net8 VSS VSS n12 l = 0.1u w = 0.96u m = 1
mmn52 nn1 SI _n5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn53 nn1 D _n7 VSS n12 l = 0.1u w = 0.21u m = 1
mmn54 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn55 net112589 NRESTORE aa VSS n12 l = 0.1u w = 0.21u m = 1
mmn56 aa jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn57 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn58 _n5 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn59 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn60 Mushegh net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn61 net155 net8 net5555555 VSS n12 l = 0.1u w = 0.21u m = 1
mmn63 net5555555 SETB net6666666 VSS n12 l = 0.1u w = 0.21u m = 1
mmn64 nn SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp30 _n8 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp31 _n6 nn VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp34 net1 VDD net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp35 net155 CLKN aa VDD p12 l = 0.1u w = 0.45u m = 1
mmp36 nn SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp37 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp38 nn1 D _n8 VDD p12 l = 0.1u w = 0.65u m = 1
mmp39 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp40 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp41 net444444 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp43 net_146 nn1 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp44 net1 net112589 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp45 net06 net_146 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp46 net112589 SETB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp47 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp48 aa jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp52 nn1 SI _n6 VDD p12 l = 0.1u w = 0.65u m = 1
mmp53 Q net8 VDD VDD p12 l = 0.1u w = 2.36u m = 1
mmp54 QN net155 VDD VDD p12 l = 0.1u w = 2.36u m = 1
mmp55 net112589 net1 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp56 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp57 net8 VDD VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp58 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp59 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp61 net155 SETB net444444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp62 net155 net8 net444444 VDD p12 l = 0.1u w = 0.33u m = 1
mmp63 net112589 RESTORE aa VDD p12 l = 0.1u w = 0.33u m = 1
mmp42 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp49 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp50 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp51 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp60 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp64 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmn38 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn43 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn46 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn48 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn50 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn62 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
.ends RSDFFSRASX2



.subckt RSDFFSRSSRX1 CLK D NRESTORE Q QN RSTB SAVE SE SETB SI VDD VDDG VSS
mmp03 net06 net0666 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp11 net2 RESTORE aa VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp19 aa jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net155 CLKN aa VDD p12 l = 0.1u w = 0.45u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp14 Q net155 VDD VDD p12 l = 0.1u w = 1.1u m = 1
mmp13 QN net8 VDD VDD p12 l = 0.1u w = 1.5u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 VDD VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp5 net1 VDD net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp12 net155 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 SET SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp16 net04 SI VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net02 RSTB net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 net05 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 net0666 net05 net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp25 net0666 SE net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 net02 D net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 net01 SET VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn03 net06 net0666 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net2 NRESTORE aa VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 VDD net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn18 aa jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKP aa VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 Q net155 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn12 net155 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 VDD net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 QN net8 VSS VSS n12 l = 0.1u w = 0.45u m = 1
mmn16 net0666 net05 net02 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 net0666 SE net04 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net04 SI VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net02 SET net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 net03 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 net02 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 SET SETB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFSRSSRX1



.subckt RSDFFSRSSRX2 CLK D NRESTORE Q QN RSTB SAVE SE SETB SI VDD VDDG VSS
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp16 net06 net05 net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp17 net04 SI VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net01 SET VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp23 net06 SE net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 net05 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp25 net02 D net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 net02 RSTB net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP n65 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 net1 VDD net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp11 net2 RESTORE _n75 VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net155 CLKN _n75 VDD p12 l = 0.1u w = 0.45u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp9 net8 VDD VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp12 net155 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 QN net8 VDD VDD p12 l = 0.1u w = 1.25u m = 2
mmp14 Q net155 VDD VDD p12 l = 0.1u w = 0.9u m = 2
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 _n75 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 SET SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp29 n65 net06 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn16 net06 SE net04 VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 net06 net05 net02 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 SET SETB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 net03 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 net04 SI VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 net02 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN n65 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 VDD net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn11 net2 NRESTORE _n75 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKP _n75 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 VDD net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net155 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 QN net8 VSS VSS n12 l = 0.1u w = 0.4u m = 2
mmn14 Q net155 VSS VSS n12 l = 0.1u w = 0.9u m = 2
mmn18 _n75 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 net02 SET net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn29 n65 net06 VSS VSS n12 l = 0.1u w = 0.21u m = 1
.ends RSDFFSRSSRX2



.subckt RSDFFSRX1 CLK D NRESTORE Q QN SAVE SE SI VDD VDDG VSS
mmp23 rrr _n53 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 0.85u m = 1
mmp12 net155 net8 net1000 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp60 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net1000 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.6u m = 1
mmp7 net155 CLKN _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp61 net1 net2 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 _n50 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 _n53 D _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5 p1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 hjf rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 p1 SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 _n53 SI net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmn24 rrr _n53 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net1 CLKN hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKP _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn60 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn61 net1 net2 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net155 net8 net1222 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.6u m = 1
mmn8 net8 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.52u m = 1
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net1222 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 _n52 p1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 _n53 SI net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n53 D _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 hjf rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 p1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFSRX1



.subckt RSDFFSRX2 CLK D NRESTORE Q QN SAVE SE SI VDD VDDG VSS
mmp23 rrr _n53 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp14 QN net155 VDD VDD p12 l = 0.1u w = 0.75u m = 2
mmp12 net155 net8 net1000 VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp60 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net1000 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp1 net1 CLKP hjf VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.6u m = 2
mmp7 net155 CLKN _n766 VDD p12 l = 0.1u w = 0.45u m = 1
mmp11 net2 RESTORE _n766 VDD p12 l = 0.1u w = 0.33u m = 1
mmp19 _n766 jk netp10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net155 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp61 net1 net2 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp18 netp10 NRESTORE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp26 RESTORE NRESTORE VDD VDD p12 l = 0.1u w = 0.48u m = 1
mmp3 _n50 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp16 _n53 D _n50 VDD p12 l = 0.1u w = 0.65u m = 1
mmp17 net5 p1 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 hjf rrr VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp24 p1 SE VDD VDD p12 l = 0.1u w = 0.55u m = 1
mmp25 _n53 SI net5 VDD p12 l = 0.1u w = 0.65u m = 1
mmn24 rrr _n53 VSS VSS n12 l = 0.1u w = 0.43u m = 1
mmn1 net1 CLKN hjf VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net155 CLKP _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn60 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn61 net1 net2 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net155 net8 net1222 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.6u m = 2
mmn8 net8 net155 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net155 VSS VSS n12 l = 0.1u w = 0.52u m = 2
mmn11 net2 NRESTORE _n766 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net1222 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn19 netn10 RESTORE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn18 _n766 jk netn10 VSS n12 l = 0.1u w = 0.21u m = 1
mmn26 RESTORE NRESTORE VSS VSS n12 l = 0.1u w = 0.24u m = 1
mmn3 _n52 p1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn16 net6 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn17 _n53 SI net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 _n53 D _n52 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 hjf rrr VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn25 p1 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 jk jk2 VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn22 SAVEN SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn21 netn102 SAVEN VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn20 jk2 jk netn102 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn32 netn103 SAVE VSS VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmn33 jk2 net8 netn103 VSS n12_hvt l = 0.1u w = 0.21u m = 1
mmp15 jk jk2 VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp22 SAVEN SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp20 netp102 SAVE VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp21 jk2 jk netp102 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp33 jk2 net8 netp103 VDDG p12_hvt l = 0.1u w = 0.33u m = 1
mmp32 netp103 SAVEN VDDG VDDG p12_hvt l = 0.1u w = 0.33u m = 1
.ends RSDFFSRX2



.subckt RSDFFX1 CLK D Q QN RETN SE SI VDD VDDG VSS
mmp26 netp26 netp22 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 netp02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp01 netp01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 INN SI netp04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp06 INP INN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 netp1 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 netp2 INP netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 INN D netp02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp6 VDD p12 l = 0.1u w = 0.41u m = 1
mmp7 netp6 CLKN VDD VDD p12 l = 0.1u w = 0.41u m = 1
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp04 netp04 netp01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 netp27 netp26 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKP netp27 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 netp5 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp103 netp103 netp102 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp105 netp102 RETN QL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp102 netp102 RETNN DL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp101 RETNN RETN VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmn26 netp26 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn06 INP INN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 netn02 netp01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 INN SI netn04 VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 netn04 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 INP netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 INN D netn02 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn6 VSS n12 l = 0.1u w = 0.23u m = 1
mmn8 netn6 CLKP VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 netp01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp27 netp26 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKN netp27 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn5 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn103 netp103 netp102 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn104 QL netp103 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn105 netp102 RETNN QL VSS n12 l = 0.1u w = 0.21u m = 1
mmn102 netp102 RETN DL VSS n12 l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends RSDFFX1



.subckt RSDFFX2 CLK D Q QN RETN SE SI VDD VDDG VSS
mmp26 netp26 netp22 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 netp02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp01 netp01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 INN SI netp04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp06 INP INN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 Q netp8 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp21 netp21 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp22 netp22 QL netp21 VDD p12 l = 0.1u w = 0.25u m = 1
mmp24 netp22 DL netp23 VDD p12 l = 0.1u w = 0.25u m = 1
mmp23 netp23 netp20 VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp1 netp1 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 netp2 INP netp1 VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 INN D netp02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 netp4 netp2 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 netp8 netp4 netp6 VDD p12 l = 0.1u w = 0.45u m = 1
mmp7 netp6 CLKN VDD VDD p12 l = 0.1u w = 0.45u m = 1
mmp9 DL netp8 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp11 QN DL VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp20 netp20 RETN VDD VDD p12 l = 0.1u w = 0.25u m = 1
mmp04 netp04 netp01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp27 netp27 netp26 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp28 netp8 CLKP netp27 VDD p12 l = 0.1u w = 0.33u m = 1
mmp5 netp5 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 netp2 netp4 netp5 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.44u m = 1
mmp103 netp103 netp102 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp104 QL netp103 VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmp105 netp102 RETN QL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp102 netp102 RETNN DL VDDG p12 l = 0.1u w = 0.33u m = 1
mmp101 RETNN RETN VDDG VDDG p12 l = 0.1u w = 0.33u m = 1
mmn26 netp26 netp22 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn06 INP INN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 netn02 netp01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 INN SI netn04 VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 netn04 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 Q netp8 VSS VSS n12 l = 0.1u w = 0.46u m = 2
mmn21 netp22 QL netn21 VSS n12 l = 0.1u w = 0.21u m = 1
mmn22 netn21 netp20 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn23 netp22 DL netn23 VSS n12 l = 0.1u w = 0.21u m = 1
mmn24 netn23 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 netn1 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 netp2 INP netn1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 netp4 netp2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 INN D netn02 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 netp8 netp4 netn6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 netn6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 DL netp8 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 QN DL VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn20 netp20 RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 netp01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn27 netp27 netp26 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn28 netp8 CLKN netp27 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 netn5 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 netp2 netp4 netn5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.22u m = 1
mmn103 netp103 netp102 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn104 QL netp103 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn105 netp102 RETNN QL VSS n12 l = 0.1u w = 0.21u m = 1
mmn102 netp102 RETN DL VSS n12 l = 0.1u w = 0.21u m = 1
mmn101 RETNN RETN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends RSDFFX2



.subckt SDFFARX1 CLK D Q QN RSTB SE SI VDD VSS
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net06 CLKP net1 VDD p12 l = 0.1u w = 0.33u m = 1
mmn1 net06 CLKN net1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.44u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.52u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1


.ends SDFFARX1



.subckt SDFFARX2 CLK D Q QN RSTB SE SI VDD VSS
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.2u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net06 CLKP net1 VDD p12 l = 0.1u w = 0.33u m = 1
mmn1 net06 CLKN net1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.76u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1


.ends SDFFARX2



.subckt SDFFASRSX1 CLK D Q QN RSTB S0 SE SETB SI VDD VSS
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp15 S0 net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.27u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 S0 net8 VSS VSS n12 l = 0.1u w = 0.45u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.45u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1


.ends SDFFASRSX1



.subckt SDFFASRSX2 CLK D Q QN RSTB S0 SE SETB SI VDD VSS
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.2u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp15 S0 net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.3u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn15 S0 net8 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1


.ends SDFFASRSX2



.subckt SDFFASRX1 CLK D Q QN RSTB SE SETB SI VDD VSS
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.27u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1


.ends SDFFASRX1



.subckt SDFFASRX2 CLK D Q QN RSTB SE SETB SI VDD VSS
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.2u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.29u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.39u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.8u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1


.ends SDFFASRX2



.subckt SDFFASX1 CLK D Q QN SE SETB SI VDD VSS
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.45u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.42u m = 1


.ends SDFFASX1



.subckt SDFFASX2 CLK D Q QN SE SETB SI VDD VSS
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.23u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.23u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.2u m = 1
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.53u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 1.12u m = 1


.ends SDFFASX2



.subckt SDFFNARX1 CLK D Q QN RSTB SE SI VDD VSS
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.5u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 0.9u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net06 CLKN net1 VDD p12 l = 0.1u w = 0.33u m = 1
mmn1 net06 CLKP net1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.35u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1


.ends SDFFNARX1



.subckt SDFFNARX2 CLK D Q QN RSTB SE SI VDD VSS
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.75u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.75u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.75u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.7u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.7u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.75u m = 1
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.75u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.7u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.75u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.75u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net06 CLKN net1 VDD p12 l = 0.1u w = 0.675u m = 1
mmn1 net06 CLKP net1 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.7u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.7u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1


.ends SDFFNARX2



.subckt SDFFNASRX1 CLK D Q QN RSTB SE SETB SI VDD VSS
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.3u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.52u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1


.ends SDFFNASRX1



.subckt SDFFNASRX2 CLK D Q QN RSTB SE SETB SI VDD VSS
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.8u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.8u m = 1
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.8u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.8u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.8u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp5 net1 RSTB net4 VDD p12 l = 0.1u w = 0.65u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.65u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.6u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp9 net8 RSTB VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.6u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.6u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKN net06 VDD p12 l = 0.1u w = 0.62u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.44u m = 1
mmn6 net1 net2 net5 VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net5 RSTB net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net8 RSTB net9 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net9 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.8u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.25u m = 1


.ends SDFFNASRX2



.subckt SDFFNASX1 CLK D Q QN SE SETB SI VDD VSS
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.6u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.45u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.6u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.5u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKN net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.4u m = 1


.ends SDFFNASX1



.subckt SDFFNASX2 CLK D Q QN SE SETB SI VDD VSS
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.61u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.65u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.65u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.65u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp3 net2 SETB VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp11 net7 SETB net10 VDD p12 l = 0.1u w = 0.65u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.65u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.59u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.3u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKN net06 VDD p12 l = 0.1u w = 0.59u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net2 SETB net3 VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net3 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net11 SETB net12 VSS n12 l = 0.1u w = 0.605u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn12 net7 net8 net11 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 1.12u m = 1


.ends SDFFNASX2



.subckt SDFFNX1 CLK D Q QN SE SI VDD VSS
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.4u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.4u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1u m = 1
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.5u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKN net06 VDD p12 l = 0.1u w = 0.5u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.33u m = 1


.ends SDFFNX1



.subckt SDFFNX2 CLK D Q QN SE SI VDD VSS
mmn10 net12 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKP net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKN net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.9u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.8u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.6u m = 1
mmp10 net10 CLKN VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.6u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.6u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.6u m = 1
mmp4 net4 CLKP VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp7 net7 CLKP net2 VDD p12 l = 0.1u w = 0.6u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKN net06 VDD p12 l = 0.1u w = 0.6u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.6u m = 1


.ends SDFFNX2



.subckt SDFFSSRX1 CLK D Q QN RSTB SE SETB SI VDD VSS
mmp05 net04 SI VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 net02 D net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 net01 SET VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net02 RSTB net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp06 net06 SE net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN IQN VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp12 IQN net8 net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp07 net05 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 IQN VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 IQN CLKN net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp08 net06 net05 net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp01 SET SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmn05 net04 SI VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net02 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 net03 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net02 SET net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn06 net06 net05 net02 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN IQN VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 IQN net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 IQN VSS VSS n12 l = 0.1u w = 0.35u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn07 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 IQN CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn08 net06 SE net04 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.5u m = 1
mmn01 SET SETB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends SDFFSSRX1



.subckt SDFFSSRX2 CLK D Q QN RSTB SE SETB SI VDD VSS
mmp05 net04 SI VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 net02 D net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp02 net01 SET VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net02 RSTB net01 VDD p12 l = 0.1u w = 0.33u m = 1
mmp06 net06 SE net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN IQN VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp12 IQN net8 net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp07 net05 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 IQN VDD VDD p12 l = 0.1u w = 0.65u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 IQN CLKN net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp08 net06 net05 net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp01 SET SETB VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmn05 net04 SI VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net02 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 net03 RSTB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net02 SET net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn06 net06 net05 net02 VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 QN IQN VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 IQN net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 IQN VSS VSS n12 l = 0.1u w = 0.35u m = 1
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn07 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 IQN CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn08 net06 SE net04 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 1u m = 1
mmn01 SET SETB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends SDFFSSRX2



.subckt SDFFX1 CLK D Q QN SE SI VDD VSS
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 0.49u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.4u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.45u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.33u m = 1


.ends SDFFX1



.subckt SDFFX2 CLK D Q QN SE SI VDD VSS
mmn10 net12 CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn8 net8 net7 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn02 net06 D net03 VSS n12 l = 0.1u w = 0.21u m = 1
mmn05 net05 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 CLKN net06 VSS n12 l = 0.1u w = 0.21u m = 1
mmn012 CLKP CLKN VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn04 net06 SI net05 VSS n12 l = 0.1u w = 0.21u m = 1
mmn03 net03 net01 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn01 net01 SE VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn011 CLKN CLK VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net1 net2 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net8 net12 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 net1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net6 CLKP VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 net7 CLKP net2 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net8 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmn14 QN net7 VSS VSS n12 l = 0.1u w = 1.12u m = 1
mmp6 net1 net2 net4 VDD p12 l = 0.1u w = 0.33u m = 1
mmp10 net10 CLKP VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp05 net06 SI net04 VDD p12 l = 0.1u w = 0.33u m = 1
mmp03 net06 D net02 VDD p12 l = 0.1u w = 0.33u m = 1
mmp12 net7 net8 net10 VDD p12 l = 0.1u w = 0.21u m = 1
mmp4 net4 CLKN VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp01 net01 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp14 QN net7 VDD VDD p12 l = 0.1u w = 2.2u m = 1
mmp011 CLKN CLK VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp2 net2 net1 VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp8 net8 net7 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp13 Q net8 VDD VDD p12 l = 0.1u w = 2.24u m = 1
mmp02 net02 SE VDD VDD p12 l = 0.1u w = 0.33u m = 1
mmp7 net7 CLKN net2 VDD p12 l = 0.1u w = 0.56u m = 1
mmp012 CLKP CLKN VDD VDD p12 l = 0.1u w = 0.21u m = 1
mmp1 net1 CLKP net06 VDD p12 l = 0.1u w = 0.33u m = 1
mmp04 net04 net01 VDD VDD p12 l = 0.1u w = 0.33u m = 1


.ends SDFFX2



.subckt SHFILL128 VDD VSS


.ends SHFILL128



.subckt SHFILL1 VDD VSS


.ends SHFILL1



.subckt SHFILL2 VDD VSS


.ends SHFILL2



.subckt SHFILL3 VDD VSS


.ends SHFILL3



.subckt SHFILL64 VDD VSS


.ends SHFILL64



.subckt TIEH VDD VSS Z
mg_pmos4t1 net1 net1 VSS VSS n12 l = 0.1u w = 0.56u m = 1
mg_nmos4t1 Z net1 VDD VDD p12 l = 0.1u w = 1.12u m = 1
.ends TIEH



.subckt TIEL VDD VSS ZN
mg_nmos4t1 net1 net1 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mg_pmos4t1 ZN net1 VSS VSS n12 l = 0.1u w = 0.56u m = 1
.ends TIEL



.subckt TNBUFFX16 ENB INP VDD VSS Z
mmn3 net3 INP VSS VSS n12 l = 0.1u w = 0.35u m = 2
mmn5 Z net3 VSS VSS n12 l = 0.1u w = 0.52u m = 16
mmn2 net2 ENB net3 VSS n12 l = 0.1u w = 0.5u m = 2
mmn4 net3 net1 VSS VSS n12 l = 0.1u w = 0.35u m = 2
mmn1 net1 ENB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 net2 INP VDD VDD p12 l = 0.1u w = 1.1u m = 2
mmp5 Z net2 VDD VDD p12 l = 0.1u w = 1.12u m = 16
mmp1 net1 ENB VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp3 net2 ENB VDD VDD p12 l = 0.1u w = 0.7u m = 2
mmp4 net3 net1 net2 VDD p12 l = 0.1u w = 0.7u m = 2


.ends TNBUFFX16



.subckt TNBUFFX1 ENB INP VDD VSS Z
mmn3 net3 INP VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn5 Z net3 VSS VSS n12 l = 0.1u w = 0.52u m = 1
mmn2 net2 ENB net3 VSS n12 l = 0.1u w = 0.35u m = 1
mmn4 net3 net1 VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn1 net1 ENB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 net2 INP VDD VDD p12 l = 0.1u w = 0.77u m = 1
mmp5 Z net2 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp1 net1 ENB VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp3 net2 ENB VDD VDD p12 l = 0.1u w = 0.49u m = 1
mmp4 net3 net1 net2 VDD p12 l = 0.1u w = 0.49u m = 1


.ends TNBUFFX1



.subckt TNBUFFX2 ENB INP VDD VSS Z
mmn3 net3 INP VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn5 Z net3 VSS VSS n12 l = 0.1u w = 0.52u m = 2
mmn2 net2 ENB net3 VSS n12 l = 0.1u w = 0.35u m = 1
mmn4 net3 net1 VSS VSS n12 l = 0.1u w = 0.25u m = 1
mmn1 net1 ENB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 net2 INP VDD VDD p12 l = 0.1u w = 0.77u m = 1
mmp5 Z net2 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp1 net1 ENB VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp3 net2 ENB VDD VDD p12 l = 0.1u w = 0.49u m = 1
mmp4 net3 net1 net2 VDD p12 l = 0.1u w = 0.49u m = 1


.ends TNBUFFX2



.subckt TNBUFFX32 ENB INP VDD VSS Z
mmn3 net3 INP VSS VSS n12 l = 0.1u w = 0.35u m = 4
mmn5 Z net3 VSS VSS n12 l = 0.1u w = 0.52u m = 32
mmn2 net2 ENB net3 VSS n12 l = 0.1u w = 0.5u m = 4
mmn4 net3 net1 VSS VSS n12 l = 0.1u w = 0.35u m = 4
mmn1 net1 ENB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 net2 INP VDD VDD p12 l = 0.1u w = 1.1u m = 4
mmp5 Z net2 VDD VDD p12 l = 0.1u w = 1.12u m = 32
mmp1 net1 ENB VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp3 net2 ENB VDD VDD p12 l = 0.1u w = 0.7u m = 4
mmp4 net3 net1 net2 VDD p12 l = 0.1u w = 0.7u m = 4


.ends TNBUFFX32



.subckt TNBUFFX4 ENB INP VDD VSS Z
mmn3 net3 INP VSS VSS n12 l = 0.1u w = 0.35u m = 1
mmn5 Z net3 VSS VSS n12 l = 0.1u w = 0.52u m = 4
mmn2 net2 ENB net3 VSS n12 l = 0.1u w = 0.5u m = 1
mmn4 net3 net1 VSS VSS n12 l = 0.1u w = 0.35u m = 1
mmn1 net1 ENB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 net2 INP VDD VDD p12 l = 0.1u w = 1.1u m = 1
mmp5 Z net2 VDD VDD p12 l = 0.1u w = 1.12u m = 4
mmp1 net1 ENB VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp3 net2 ENB VDD VDD p12 l = 0.1u w = 0.7u m = 1
mmp4 net3 net1 net2 VDD p12 l = 0.1u w = 0.7u m = 1


.ends TNBUFFX4



.subckt TNBUFFX8 ENB INP VDD VSS Z
mmn3 net3 INP VSS VSS n12 l = 0.1u w = 0.35u m = 1
mmn5 Z net3 VSS VSS n12 l = 0.1u w = 0.52u m = 8
mmn2 net2 ENB net3 VSS n12 l = 0.1u w = 0.5u m = 1
mmn4 net3 net1 VSS VSS n12 l = 0.1u w = 0.35u m = 1
mmn1 net1 ENB VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmp2 net2 INP VDD VDD p12 l = 0.1u w = 1.1u m = 1
mmp5 Z net2 VDD VDD p12 l = 0.1u w = 1.12u m = 8
mmp1 net1 ENB VDD VDD p12 l = 0.1u w = 0.5u m = 1
mmp3 net2 ENB VDD VDD p12 l = 0.1u w = 0.7u m = 1
mmp4 net3 net1 net2 VDD p12 l = 0.1u w = 0.7u m = 1


.ends TNBUFFX8



.subckt XOR3X2_LVT 
M_MMN2 NET2 IN2 VSS VSS n12_lvt  l=0.100u w=0.230u
M_MMN7 NET7 IN3 VSS VSS n12_lvt  l=0.100u w=0.210u
M_ld_M3 VSS NET11 Q VSS n12_lvt  l=0.100u w=0.490u
M_ld_M4 Q NET11 VSS VSS n12_lvt  l=0.100u w=0.490u
M_MMN8 VSS NET8 NET9 VSS n12_lvt  l=0.100u w=0.140u
M_ld_M6 NET4 NET1 NET8 VSS n12_lvt  l=0.100u w=0.230u
M_ld_M7 NET4 NET2 VSS VSS n12_lvt  l=0.100u w=0.230u
M_ld_M8 VSS IN2 NET6 VSS n12_lvt  l=0.100u w=0.230u
M_MMN1 VSS IN1 NET1 VSS n12_lvt  l=0.100u w=0.230u
M_ld_M10 NET8 IN1 NET6 VSS n12_lvt  l=0.100u w=0.230u
M_MMN10 NET8 IN3 NET11 VSS n12_lvt  l=0.100u w=0.140u
M_MMN9 NET9 NET7 NET11 VSS n12_lvt  l=0.100u w=0.140u
M_MMP10 NET11 NET7 NET8 VDD p12_lvt  l=0.100u w=0.580u
M_MMP9 NET11 IN3 NET9 VDD p12_lvt  l=0.100u w=0.580u
M_MMP2 NET2 IN2 VDD VDD p12_lvt  l=0.100u w=0.420u
M_MMP7 NET7 IN3 VDD VDD p12_lvt  l=0.100u w=0.350u
M_MMP8 NET9 NET8 VDD VDD p12_lvt  l=0.100u w=0.350u
M_MMP1 NET1 IN1 VDD VDD p12_lvt  l=0.100u w=0.420u
M_ld_M19 VDD NET11 Q VDD p12_lvt  l=0.100u w=1.120u
M_ld_M20 Q NET11 VDD VDD p12_lvt  l=0.100u w=1.120u
M_ld_M21 NET3 NET1 NET8 VDD p12_lvt  l=0.100u w=0.640u
M_ld_M22 VDD NET2 NET5 VDD p12_lvt  l=0.100u w=0.640u
M_ld_M23 NET3 IN2 VDD VDD p12_lvt  l=0.100u w=0.640u
M_ld_M24 NET8 IN1 NET5 VDD p12_lvt  l=0.100u w=0.640u
.ends XOR3X2_LVT

.subckt XNOR2X1 IN1 IN2 Q VDD VSS
mmp4 net7 net1 net3 VDD p12 l = 0.1u w = 0.6u m = 1
mmp5 net5 net2 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp3 net3 IN2 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp6 net7 IN1 net5 VDD p12 l = 0.1u w = 0.6u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.32u m = 1
mmp7 Q net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp2 net2 IN2 VDD VDD p12 l = 0.1u w = 0.32u m = 1
mmn3 net7 net1 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net4 net2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 Q net7 VSS VSS n12 l = 0.1u w = 0.42u m = 1
mmn1 net1 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net6 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net7 IN1 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends XNOR2X1



.subckt XNOR2X2 IN1 IN2 Q VDD VSS
mmp8 net2 IN2 VDD VDD p12 l = 0.1u w = 0.32u m = 1
mmp9 net5 net2 VDD VDD p12 l = 0.1u w = 0.62u m = 1
mmp10 net7 IN1 net5 VDD p12 l = 0.1u w = 0.62u m = 1
mmp11 net1 IN1 VDD VDD p12 l = 0.1u w = 0.32u m = 1
mmp12 net7 net1 net3 VDD p12 l = 0.1u w = 0.62u m = 1
mmp13 net3 IN2 VDD VDD p12 l = 0.1u w = 0.62u m = 1
mmp14 Q net7 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmn8 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn9 net6 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net4 net2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net7 IN1 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net7 net1 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 Q net7 VSS VSS n12 l = 0.1u w = 0.42u m = 2
mmn14 net1 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1


.ends XNOR2X2



.subckt XNOR3X1 IN1 IN2 IN3 Q VDD VSS
mmn10 net10 IN3 net11 VSS n12 l = 0.1u w = 0.14u m = 1
mmn3 net8 net1 net4 VSS n12 l = 0.1u w = 0.23u m = 1
mmn9 net8 net7 net11 VSS n12 l = 0.1u w = 0.14u m = 1
mmn11 Q net11 VSS VSS n12 l = 0.1u w = 0.44u m = 1
mmn7 net7 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn5 net8 IN1 net6 VSS n12 l = 0.1u w = 0.23u m = 1
mmn6 net6 IN2 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn1 net1 IN1 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn8 net10 net8 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn4 net4 net2 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmp9 net8 IN3 net11 VDD p12 l = 0.1u w = 0.52u m = 1
mmp3 net3 IN2 VDD VDD p12 l = 0.1u w = 0.64u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp5 net5 net2 VDD VDD p12 l = 0.1u w = 0.64u m = 1
mmp10 net10 net7 net11 VDD p12 l = 0.1u w = 0.52u m = 1
mmp4 net8 net1 net3 VDD p12 l = 0.1u w = 0.64u m = 1
mmp7 net7 IN3 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp8 net10 net8 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp11 Q net11 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmp6 net8 IN1 net5 VDD p12 l = 0.1u w = 0.64u m = 1
mmp2 net2 IN2 VDD VDD p12 l = 0.1u w = 0.42u m = 1


.ends XNOR3X1



.subckt XNOR3X2 IN1 IN2 IN3 Q VDD VSS
mmp2 net2 IN2 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp8 net10 net8 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp3 net3 IN2 VDD VDD p12 l = 0.1u w = 0.64u m = 1
mmp10 net10 net7 net11 VDD p12 l = 0.1u w = 0.58u m = 1
mmp7 net7 IN3 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp4 net8 net1 net3 VDD p12 l = 0.1u w = 0.64u m = 1
mmp6 net8 IN1 net5 VDD p12 l = 0.1u w = 0.64u m = 1
mmp5 net5 net2 VDD VDD p12 l = 0.1u w = 0.64u m = 1
mmp11 Q net11 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp9 net8 IN3 net11 VDD p12 l = 0.1u w = 0.58u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmn9 net8 net7 net11 VSS n12 l = 0.1u w = 0.14u m = 1
mmn3 net8 net1 net4 VSS n12 l = 0.1u w = 0.23u m = 1
mmn8 net10 net8 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn5 net8 IN1 net6 VSS n12 l = 0.1u w = 0.23u m = 1
mmn7 net7 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 IN1 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn4 net4 net2 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn10 net10 IN3 net11 VSS n12 l = 0.1u w = 0.14u m = 1
mmn11 Q net11 VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn6 net6 IN2 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.23u m = 1


.ends XNOR3X2



.subckt XOR2X1 IN1 IN2 Q VDD VSS
mmp2 net2 IN2 VDD VDD p12 l = 0.1u w = 0.32u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.32u m = 1
mmp3 net3 IN2 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp4 net7 IN1 net3 VDD p12 l = 0.1u w = 0.6u m = 1
mmp5 net5 net2 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp6 net7 net1 net5 VDD p12 l = 0.1u w = 0.6u m = 1
mmp7 Q net7 VDD VDD p12 l = 0.1u w = 1.12u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net7 IN1 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn1 net1 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn4 net4 net2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn5 net7 net1 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmn6 net6 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn7 Q net7 VSS VSS n12 l = 0.1u w = 0.4u m = 1


.ends XOR2X1



.subckt XOR2X2 IN1 IN2 Q VDD VSS
mmn8 Q net7 VSS VSS n12 l = 0.1u w = 0.4u m = 2
mmn9 net6 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn10 net7 IN1 net4 VSS n12 l = 0.1u w = 0.21u m = 1
mmn11 net1 IN1 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn12 net4 net2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn13 net2 IN2 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 net7 net1 net6 VSS n12 l = 0.1u w = 0.21u m = 1
mmp8 net7 IN1 net3 VDD p12 l = 0.1u w = 0.6u m = 1
mmp9 Q net7 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp10 net2 IN2 VDD VDD p12 l = 0.1u w = 0.32u m = 1
mmp11 net3 IN2 VDD VDD p12 l = 0.1u w = 0.6u m = 1
mmp12 net7 net1 net5 VDD p12 l = 0.1u w = 0.6u m = 1
mmp13 net1 IN1 VDD VDD p12 l = 0.1u w = 0.32u m = 1
mmp14 net5 net2 VDD VDD p12 l = 0.1u w = 0.6u m = 1


.ends XOR2X2



.subckt XOR3X1 IN1 IN2 IN3 Q VDD VSS
mmn6 net6 IN2 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn7 net7 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn3 net8 net1 net4 VSS n12 l = 0.1u w = 0.23u m = 1
mmn4 net4 net2 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn5 net8 IN1 net6 VSS n12 l = 0.1u w = 0.23u m = 1
mmn2 net2 IN2 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn1 net1 IN1 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn9 net9 net7 net11 VSS n12 l = 0.1u w = 0.14u m = 1
mmn10 net8 IN3 net11 VSS n12 l = 0.1u w = 0.14u m = 1
mmn8 net9 net8 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn11 Q net11 VSS VSS n12 l = 0.1u w = 0.44u m = 1
mmp1 net1 IN1 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp4 net8 net1 net3 VDD p12 l = 0.1u w = 0.64u m = 1
mmp2 net2 IN2 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp6 net8 IN1 net5 VDD p12 l = 0.1u w = 0.64u m = 1
mmp3 net3 IN2 VDD VDD p12 l = 0.1u w = 0.64u m = 1
mmp7 net7 IN3 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp5 net5 net2 VDD VDD p12 l = 0.1u w = 0.64u m = 1
mmp9 net9 IN3 net11 VDD p12 l = 0.1u w = 0.52u m = 1
mmp10 net8 net7 net11 VDD p12 l = 0.1u w = 0.52u m = 1
mmp8 net9 net8 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp11 Q net11 VDD VDD p12 l = 0.1u w = 1.12u m = 1


.ends XOR3X1



.subckt XOR3X2 IN1 IN2 IN3 Q VDD VSS
mmn12 net4 net2 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn13 net7 IN3 VSS VSS n12 l = 0.1u w = 0.21u m = 1
mmn14 net2 IN2 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn15 net8 net1 net4 VSS n12 l = 0.1u w = 0.23u m = 1
mmn16 net9 net8 VSS VSS n12 l = 0.1u w = 0.14u m = 1
mmn17 net8 IN3 net11 VSS n12 l = 0.1u w = 0.14u m = 1
mmn18 net8 IN1 net6 VSS n12 l = 0.1u w = 0.23u m = 1
mmn19 net9 net7 net11 VSS n12 l = 0.1u w = 0.14u m = 1
mmn20 Q net11 VSS VSS n12 l = 0.1u w = 0.5u m = 2
mmn21 net1 IN1 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmn22 net6 IN2 VSS VSS n12 l = 0.1u w = 0.23u m = 1
mmp12 net8 net7 net11 VDD p12 l = 0.1u w = 0.58u m = 1
mmp13 net7 IN3 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp14 net5 net2 VDD VDD p12 l = 0.1u w = 0.64u m = 1
mmp15 net1 IN1 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp16 net9 net8 VDD VDD p12 l = 0.1u w = 0.35u m = 1
mmp17 net8 net1 net3 VDD p12 l = 0.1u w = 0.64u m = 1
mmp18 net8 IN1 net5 VDD p12 l = 0.1u w = 0.64u m = 1
mmp19 net2 IN2 VDD VDD p12 l = 0.1u w = 0.42u m = 1
mmp20 Q net11 VDD VDD p12 l = 0.1u w = 1.12u m = 2
mmp21 net3 IN2 VDD VDD p12 l = 0.1u w = 0.64u m = 1
mmp22 net9 IN3 net11 VDD p12 l = 0.1u w = 0.58u m = 1


.ends XOR3X2


