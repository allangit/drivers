
module multi_reloj_N_filtros8 (filtro_pipelining_clk_2x , reset , 
    reloj_secuencia );
input  filtro_pipelining_clk_2x ;
input  reset ;
output [7:0] reloj_secuencia ;


wire [7:2] add_x_58_1_carry ;

DFFARX1 contador_reg_2_ (.CLK ( filtro_pipelining_clk_2x ) , .RSTB ( n8 ) 
    , .QN ( n6 ) , .Q ( reloj_secuencia[2] ) , .D ( N3 ) ) ;
DFFARX1 contador_reg_3_ (.CLK ( filtro_pipelining_clk_2x ) , .RSTB ( n8 ) 
    , .QN ( n3 ) , .Q ( reloj_secuencia[3] ) , .D ( N4 ) ) ;
DFFARX1 contador_reg_4_ (.CLK ( filtro_pipelining_clk_2x ) , .RSTB ( n8 ) 
    , .QN ( n5 ) , .Q ( reloj_secuencia[4] ) , .D ( N5 ) ) ;
DFFARX1 contador_reg_5_ (.CLK ( filtro_pipelining_clk_2x ) , .RSTB ( n8 ) 
    , .QN ( n4 ) , .Q ( reloj_secuencia[5] ) , .D ( N6 ) ) ;
DFFARX1 contador_reg_6_ (.CLK ( filtro_pipelining_clk_2x ) , .RSTB ( n8 ) 
    , .QN ( n2 ) , .Q ( reloj_secuencia[6] ) , .D ( N7 ) ) ;
DFFARX1 contador_reg_7_ (.CLK ( filtro_pipelining_clk_2x ) , .RSTB ( n8 ) 
    , .QN ( n1 ) , .Q ( reloj_secuencia[7] ) , .D ( N8 ) ) ;
INVX0 U3 (.ZN ( n8 ) , .INP ( reset ) ) ;
HADDX1 add_x_58_1_U1_1_6 (.B0 ( add_x_58_1_carry[6] ) 
    , .A0 ( add_x_58_1_A_6_ ) , .C1 ( add_x_58_1_carry[7] ) , .SO ( N7 ) ) ;
HADDX1 add_x_58_1_U1_1_5 (.B0 ( add_x_58_1_carry[5] ) 
    , .A0 ( add_x_58_1_A_5_ ) , .C1 ( add_x_58_1_carry[6] ) , .SO ( N6 ) ) ;
HADDX1 add_x_58_1_U1_1_4 (.B0 ( add_x_58_1_carry[4] ) 
    , .A0 ( add_x_58_1_A_4_ ) , .C1 ( add_x_58_1_carry[5] ) , .SO ( N5 ) ) ;
HADDX1 add_x_58_1_U1_1_3 (.B0 ( add_x_58_1_carry[3] ) 
    , .A0 ( add_x_58_1_A_3_ ) , .C1 ( add_x_58_1_carry[4] ) , .SO ( N4 ) ) ;
HADDX1 add_x_58_1_U1_1_2 (.B0 ( add_x_58_1_carry[2] ) 
    , .A0 ( add_x_58_1_A_2_ ) , .C1 ( add_x_58_1_carry[3] ) , .SO ( N3 ) ) ;
DFFARX1 contador_reg_0_ (.CLK ( filtro_pipelining_clk_2x ) , .RSTB ( n8 ) 
    , .QN ( n7 ) , .Q ( reloj_secuencia[0] ) , .D ( n7 ) ) ;
DFFARX1 contador_reg_1_ (.CLK ( filtro_pipelining_clk_2x ) , .RSTB ( n8 ) 
    , .QN ( n9 ) , .Q ( reloj_secuencia[1] ) , .D ( N2 ) ) ;
INVX0 U11 (.ZN ( add_x_58_1_A_2_ ) , .INP ( n6 ) ) ;
INVX0 U10 (.ZN ( add_x_58_1_A_4_ ) , .INP ( n5 ) ) ;
INVX0 U9 (.ZN ( add_x_58_1_A_5_ ) , .INP ( n4 ) ) ;
INVX0 U8 (.ZN ( add_x_58_1_A_3_ ) , .INP ( n3 ) ) ;
INVX0 U7 (.ZN ( add_x_58_1_A_6_ ) , .INP ( n2 ) ) ;
XNOR2X1 U6 (.IN1 ( n1 ) , .IN2 ( add_x_58_1_carry[7] ) , .Q ( N8 ) ) ;
NOR2X0 U5 (.QN ( add_x_58_1_carry[2] ) , .IN1 ( n7 ) , .IN2 ( n9 ) ) ;
XOR2X1 U4 (.IN2 ( n9 ) , .Q ( N2 ) , .IN1 ( n7 ) ) ;
endmodule




module filtro_pipelining (filtro_pipelining_in , filtro_pipelining_salida , 
    reset , filtro_pipelining_clk_2x );
input  [15:0] filtro_pipelining_in ;
output [127:0] filtro_pipelining_salida ;
input  reset ;
input  filtro_pipelining_clk_2x ;

wire [7:0] reloj_secuencia ;

wire [141:0] bank_registro_registros ;
wire [18:0] partial_1 ;
wire [18:0] sos2_reg_entrada ;
wire [6:0] reloj_secuencia_delay ;
wire [18:0] bajo_reg_entrada ;
wire [15:0] alto_reg_entrada ;
wire [18:0] partial_2_L ;
wire [18:0] partial_2_H ;
wire [18:2] partial_3_H ;
wire [18:2] partial_3_L ;
wire [17:0] coeficiente_b12_H_v_out ;
wire [17:0] coeficiente_b12_L_v_out ;
wire [17:0] in_reg_salida_v ;
wire [18:0] coeficiente_a22_in ;
wire [18:0] coeficiente_b11_H_v_out ;
wire [18:0] coeficiente_b11_L_v_out ;
wire [18:10] coeficiente_a11_H_in ;


multi_reloj_N_filtros8 multi_reloj (
    .filtro_pipelining_clk_2x ( filtro_pipelining_clk_2x ) , .reset ( reset ) , 
    .reloj_secuencia ( reloj_secuencia ) ) ;

DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1657 ) 
    , .Q ( bank_registro_registros[3] ) , .D ( filtro_pipelining_in[3] ) ) ;
DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1656 ) 
    , .Q ( bank_registro_registros[2] ) , .D ( filtro_pipelining_in[2] ) ) ;
DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1646 ) 
    , .Q ( bank_registro_registros[1] ) , .D ( filtro_pipelining_in[1] ) ) ;
DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1659 ) 
    , .Q ( bank_registro_registros[0] ) , .D ( filtro_pipelining_in[0] ) ) ;
DFFNX1 secuencia_reloj_prioridad_salida_reg_1_ (
    .CLK ( filtro_pipelining_clk_2x ) 
    , .D ( secuencia_reloj_prioridad_salida_pre_1_ ) , .QN ( n1491 ) 
    , .Q ( seleccion_1_ ) ) ;
DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1657 ) 
    , .Q ( bank_registro_registros[11] ) , .D ( filtro_pipelining_in[11] ) ) ;
DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1656 ) 
    , .Q ( bank_registro_registros[10] ) , .D ( filtro_pipelining_in[10] ) ) ;
DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1654 ) 
    , .Q ( bank_registro_registros[9] ) , .D ( filtro_pipelining_in[9] ) ) ;
DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1655 ) 
    , .Q ( bank_registro_registros[8] ) , .D ( filtro_pipelining_in[8] ) ) ;
DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1657 ) 
    , .Q ( bank_registro_registros[7] ) , .D ( filtro_pipelining_in[7] ) ) ;
DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1656 ) 
    , .Q ( bank_registro_registros[6] ) , .D ( filtro_pipelining_in[6] ) ) ;
DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1654 ) 
    , .Q ( bank_registro_registros[5] ) , .D ( filtro_pipelining_in[5] ) ) ;
DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1655 ) 
    , .Q ( bank_registro_registros[4] ) , .D ( filtro_pipelining_in[4] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][3] ) , .D ( partial_1[3] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][2] ) , .D ( partial_1[2] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][1] ) , .D ( partial_1[1] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][0] ) , .D ( partial_1[0] ) ) ;
DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1654 ) 
    , .Q ( bank_registro_registros[15] ) , .D ( filtro_pipelining_in[15] ) ) ;
DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1657 ) 
    , .Q ( bank_registro_registros[14] ) , .D ( filtro_pipelining_in[14] ) ) ;
DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1655 ) 
    , .Q ( bank_registro_registros[13] ) , .D ( filtro_pipelining_in[13] ) ) ;
DFFARX1 in_reg_pila_registro_reg_0_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1655 ) 
    , .Q ( bank_registro_registros[12] ) , .D ( filtro_pipelining_in[12] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][11] ) , .D ( partial_1[11] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][10] ) , .D ( partial_1[10] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][9] ) , .D ( partial_1[9] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][8] ) , .D ( partial_1[8] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][7] ) , .D ( partial_1[7] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][6] ) , .D ( partial_1[6] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][5] ) , .D ( partial_1[5] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][4] ) , .D ( partial_1[4] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][0] ) , .D ( partial_1[0] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][18] ) , .D ( partial_1[18] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][17] ) , .D ( partial_1[17] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][16] ) , .D ( partial_1[16] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][15] ) , .D ( partial_1[15] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][14] ) , .D ( partial_1[14] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][13] ) , .D ( partial_1[13] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_0_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[0][12] ) , .D ( partial_1[12] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][8] ) , .D ( partial_1[8] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][7] ) , .D ( partial_1[7] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][6] ) , .D ( partial_1[6] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][5] ) , .D ( partial_1[5] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][4] ) , .D ( partial_1[4] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][3] ) , .D ( partial_1[3] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][2] ) , .D ( partial_1[2] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][1] ) , .D ( partial_1[1] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][16] ) , .D ( partial_1[16] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][15] ) , .D ( partial_1[15] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][14] ) , .D ( partial_1[14] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][13] ) , .D ( partial_1[13] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][12] ) , .D ( partial_1[12] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][11] ) , .D ( partial_1[11] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][10] ) , .D ( partial_1[10] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][9] ) , .D ( partial_1[9] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][5] ) , .D ( partial_1[5] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][4] ) , .D ( partial_1[4] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][3] ) , .D ( partial_1[3] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][2] ) , .D ( partial_1[2] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][1] ) , .D ( partial_1[1] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][0] ) , .D ( partial_1[0] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][18] ) , .D ( partial_1[18] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_1_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[1][17] ) , .D ( partial_1[17] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][13] ) , .D ( partial_1[13] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][12] ) , .D ( partial_1[12] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][11] ) , .D ( partial_1[11] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][10] ) , .D ( partial_1[10] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][9] ) , .D ( partial_1[9] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][8] ) , .D ( partial_1[8] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][7] ) , .D ( partial_1[7] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][6] ) , .D ( partial_1[6] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][2] ) , .D ( partial_1[2] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][1] ) , .D ( partial_1[1] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][0] ) , .D ( partial_1[0] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][18] ) , .D ( partial_1[18] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][17] ) , .D ( partial_1[17] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][16] ) , .D ( partial_1[16] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][15] ) , .D ( partial_1[15] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_2_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[2][14] ) , .D ( partial_1[14] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][10] ) , .D ( partial_1[10] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][9] ) , .D ( partial_1[9] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][8] ) , .D ( partial_1[8] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][7] ) , .D ( partial_1[7] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][6] ) , .D ( partial_1[6] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][5] ) , .D ( partial_1[5] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][4] ) , .D ( partial_1[4] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][3] ) , .D ( partial_1[3] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][18] ) , .D ( partial_1[18] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][17] ) , .D ( partial_1[17] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][16] ) , .D ( partial_1[16] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][15] ) , .D ( partial_1[15] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][14] ) , .D ( partial_1[14] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][13] ) , .D ( partial_1[13] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][12] ) , .D ( partial_1[12] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_3_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[3][11] ) , .D ( partial_1[11] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][7] ) , .D ( partial_1[7] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][6] ) , .D ( partial_1[6] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][5] ) , .D ( partial_1[5] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][4] ) , .D ( partial_1[4] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][3] ) , .D ( partial_1[3] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][2] ) , .D ( partial_1[2] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][1] ) , .D ( partial_1[1] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][0] ) , .D ( partial_1[0] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][15] ) , .D ( partial_1[15] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][14] ) , .D ( partial_1[14] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][13] ) , .D ( partial_1[13] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][12] ) , .D ( partial_1[12] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][11] ) , .D ( partial_1[11] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][10] ) , .D ( partial_1[10] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][9] ) , .D ( partial_1[9] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1654 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][8] ) , .D ( partial_1[8] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][4] ) , .D ( partial_1[4] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][3] ) , .D ( partial_1[3] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][2] ) , .D ( partial_1[2] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][1] ) , .D ( partial_1[1] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][0] ) , .D ( partial_1[0] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][18] ) , .D ( partial_1[18] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][17] ) , .D ( partial_1[17] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_4_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[4][16] ) , .D ( partial_1[16] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][12] ) , .D ( partial_1[12] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][11] ) , .D ( partial_1[11] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][10] ) , .D ( partial_1[10] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][9] ) , .D ( partial_1[9] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][8] ) , .D ( partial_1[8] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][7] ) , .D ( partial_1[7] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][6] ) , .D ( partial_1[6] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][5] ) , .D ( partial_1[5] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][1] ) , .D ( partial_1[1] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][0] ) , .D ( partial_1[0] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][18] ) , .D ( partial_1[18] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][17] ) , .D ( partial_1[17] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][16] ) , .D ( partial_1[16] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][15] ) , .D ( partial_1[15] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][14] ) , .D ( partial_1[14] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_5_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[5][13] ) , .D ( partial_1[13] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][9] ) , .D ( partial_1[9] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][8] ) , .D ( partial_1[8] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][7] ) , .D ( partial_1[7] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][6] ) , .D ( partial_1[6] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][5] ) , .D ( partial_1[5] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][4] ) , .D ( partial_1[4] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][3] ) , .D ( partial_1[3] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][2] ) , .D ( partial_1[2] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][17] ) , .D ( partial_1[17] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][16] ) , .D ( partial_1[16] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][15] ) , .D ( partial_1[15] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][14] ) , .D ( partial_1[14] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][13] ) , .D ( partial_1[13] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][12] ) , .D ( partial_1[12] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][11] ) , .D ( partial_1[11] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][10] ) , .D ( partial_1[10] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1659 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][1] ) , .D ( sos2_reg_entrada[1] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1659 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][1] ) , .D ( sos2_reg_entrada[1] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1658 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][1] ) , .D ( sos2_reg_entrada[1] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1658 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][1] ) , .D ( sos2_reg_entrada[1] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][1] ) , .D ( partial_1[1] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1659 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][0] ) , .D ( sos2_reg_entrada[0] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1658 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][0] ) , .D ( partial_1[0] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_6_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1659 ) 
    , .Q ( \sos1_reg/bank_registro_registros[6][18] ) , .D ( partial_1[18] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1657 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][2] ) , .D ( sos2_reg_entrada[2] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1656 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][2] ) , .D ( sos2_reg_entrada[2] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][2] ) , .D ( sos2_reg_entrada[2] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][2] ) , .D ( partial_1[2] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1656 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][1] ) , .D ( sos2_reg_entrada[1] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][1] ) , .D ( sos2_reg_entrada[1] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1655 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][1] ) , .D ( sos2_reg_entrada[1] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1657 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][1] ) , .D ( sos2_reg_entrada[1] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1655 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][3] ) , .D ( sos2_reg_entrada[3] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][3] ) , .D ( sos2_reg_entrada[3] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][3] ) , .D ( partial_1[3] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1657 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][2] ) , .D ( sos2_reg_entrada[2] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1655 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][2] ) , .D ( sos2_reg_entrada[2] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1656 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][2] ) , .D ( sos2_reg_entrada[2] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][2] ) , .D ( sos2_reg_entrada[2] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1655 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][2] ) , .D ( sos2_reg_entrada[2] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1656 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][4] ) , .D ( sos2_reg_entrada[4] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][4] ) , .D ( partial_1[4] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1656 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][3] ) , .D ( sos2_reg_entrada[3] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][3] ) , .D ( sos2_reg_entrada[3] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][3] ) , .D ( sos2_reg_entrada[3] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1655 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][3] ) , .D ( sos2_reg_entrada[3] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1656 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][3] ) , .D ( sos2_reg_entrada[3] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1657 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][3] ) , .D ( sos2_reg_entrada[3] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1655 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][5] ) , .D ( partial_1[5] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][4] ) , .D ( sos2_reg_entrada[4] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1655 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][4] ) , .D ( sos2_reg_entrada[4] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1657 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][4] ) , .D ( sos2_reg_entrada[4] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1656 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][4] ) , .D ( sos2_reg_entrada[4] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1655 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][4] ) , .D ( sos2_reg_entrada[4] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1657 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][4] ) , .D ( sos2_reg_entrada[4] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][4] ) , .D ( sos2_reg_entrada[4] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1656 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][5] ) , .D ( sos2_reg_entrada[5] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][5] ) , .D ( sos2_reg_entrada[5] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1655 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][5] ) , .D ( sos2_reg_entrada[5] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1657 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][5] ) , .D ( sos2_reg_entrada[5] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1656 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][5] ) , .D ( sos2_reg_entrada[5] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1656 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][5] ) , .D ( sos2_reg_entrada[5] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][5] ) , .D ( sos2_reg_entrada[5] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][5] ) , .D ( sos2_reg_entrada[5] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1655 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][6] ) , .D ( sos2_reg_entrada[6] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][6] ) , .D ( sos2_reg_entrada[6] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1655 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][6] ) , .D ( sos2_reg_entrada[6] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1657 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][6] ) , .D ( sos2_reg_entrada[6] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1656 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][6] ) , .D ( sos2_reg_entrada[6] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][6] ) , .D ( sos2_reg_entrada[6] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1655 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][6] ) , .D ( sos2_reg_entrada[6] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][6] ) , .D ( partial_1[6] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1655 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][7] ) , .D ( sos2_reg_entrada[7] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1657 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][7] ) , .D ( sos2_reg_entrada[7] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1656 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][7] ) , .D ( sos2_reg_entrada[7] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][7] ) , .D ( sos2_reg_entrada[7] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1655 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][7] ) , .D ( sos2_reg_entrada[7] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1657 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][7] ) , .D ( sos2_reg_entrada[7] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1656 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][7] ) , .D ( partial_1[7] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][6] ) , .D ( sos2_reg_entrada[6] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1649 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][8] ) , .D ( sos2_reg_entrada[8] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1649 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][8] ) , .D ( sos2_reg_entrada[8] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1649 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][8] ) , .D ( sos2_reg_entrada[8] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1655 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][8] ) , .D ( sos2_reg_entrada[8] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][8] ) , .D ( sos2_reg_entrada[8] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1657 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][8] ) , .D ( partial_1[8] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1656 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][7] ) , .D ( sos2_reg_entrada[7] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1654 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][7] ) , .D ( sos2_reg_entrada[7] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][9] ) , .D ( sos2_reg_entrada[9] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][9] ) , .D ( sos2_reg_entrada[9] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][9] ) , .D ( sos2_reg_entrada[9] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][9] ) , .D ( sos2_reg_entrada[9] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1648 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][9] ) , .D ( partial_1[9] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][8] ) , .D ( sos2_reg_entrada[8] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][8] ) , .D ( sos2_reg_entrada[8] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1649 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][8] ) , .D ( sos2_reg_entrada[8] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1651 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][10] ) 
    , .D ( sos2_reg_entrada[10] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1650 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][10] ) 
    , .D ( sos2_reg_entrada[10] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1649 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][10] ) 
    , .D ( sos2_reg_entrada[10] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1648 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][10] ) , .D ( partial_1[10] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][9] ) , .D ( sos2_reg_entrada[9] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][9] ) , .D ( sos2_reg_entrada[9] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][9] ) , .D ( sos2_reg_entrada[9] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][9] ) , .D ( sos2_reg_entrada[9] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1653 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][11] ) 
    , .D ( sos2_reg_entrada[11] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1651 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][11] ) 
    , .D ( sos2_reg_entrada[11] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1650 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][11] ) , .D ( partial_1[11] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1649 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][10] ) 
    , .D ( sos2_reg_entrada[10] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][10] ) 
    , .D ( sos2_reg_entrada[10] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1652 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][10] ) 
    , .D ( sos2_reg_entrada[10] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1647 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][10] ) 
    , .D ( sos2_reg_entrada[10] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1653 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][10] ) 
    , .D ( sos2_reg_entrada[10] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][12] ) 
    , .D ( sos2_reg_entrada[12] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1648 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][12] ) , .D ( partial_1[12] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][11] ) 
    , .D ( sos2_reg_entrada[11] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][11] ) 
    , .D ( sos2_reg_entrada[11] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][11] ) 
    , .D ( sos2_reg_entrada[11] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][11] ) 
    , .D ( sos2_reg_entrada[11] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][11] ) 
    , .D ( sos2_reg_entrada[11] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1647 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][11] ) 
    , .D ( sos2_reg_entrada[11] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1661 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][13] ) , .D ( partial_1[13] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1651 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][12] ) 
    , .D ( sos2_reg_entrada[12] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1663 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][12] ) 
    , .D ( sos2_reg_entrada[12] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][12] ) 
    , .D ( sos2_reg_entrada[12] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][12] ) 
    , .D ( sos2_reg_entrada[12] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][12] ) 
    , .D ( sos2_reg_entrada[12] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][12] ) 
    , .D ( sos2_reg_entrada[12] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][12] ) 
    , .D ( sos2_reg_entrada[12] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1660 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][13] ) 
    , .D ( sos2_reg_entrada[13] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1659 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][13] ) 
    , .D ( sos2_reg_entrada[13] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1650 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][13] ) 
    , .D ( sos2_reg_entrada[13] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1647 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][13] ) 
    , .D ( sos2_reg_entrada[13] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1658 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][13] ) 
    , .D ( sos2_reg_entrada[13] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1659 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][13] ) 
    , .D ( sos2_reg_entrada[13] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1649 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][13] ) 
    , .D ( sos2_reg_entrada[13] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1653 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][13] ) 
    , .D ( sos2_reg_entrada[13] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][14] ) 
    , .D ( sos2_reg_entrada[14] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][14] ) 
    , .D ( sos2_reg_entrada[14] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][14] ) 
    , .D ( sos2_reg_entrada[14] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][14] ) 
    , .D ( sos2_reg_entrada[14] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][14] ) 
    , .D ( sos2_reg_entrada[14] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][14] ) 
    , .D ( sos2_reg_entrada[14] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][14] ) 
    , .D ( sos2_reg_entrada[14] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1662 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][14] ) , .D ( partial_1[14] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1647 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][15] ) 
    , .D ( sos2_reg_entrada[15] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1647 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][15] ) 
    , .D ( sos2_reg_entrada[15] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1647 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][15] ) 
    , .D ( sos2_reg_entrada[15] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1647 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][15] ) 
    , .D ( sos2_reg_entrada[15] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][15] ) 
    , .D ( sos2_reg_entrada[15] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][15] ) 
    , .D ( sos2_reg_entrada[15] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1648 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][15] ) , .D ( partial_1[15] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][14] ) 
    , .D ( sos2_reg_entrada[14] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1647 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][16] ) 
    , .D ( sos2_reg_entrada[16] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1647 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][16] ) 
    , .D ( sos2_reg_entrada[16] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1647 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][16] ) 
    , .D ( sos2_reg_entrada[16] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1647 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][16] ) 
    , .D ( sos2_reg_entrada[16] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1647 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][16] ) 
    , .D ( sos2_reg_entrada[16] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1647 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][16] ) , .D ( partial_1[16] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1647 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][15] ) 
    , .D ( sos2_reg_entrada[15] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1647 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][15] ) 
    , .D ( sos2_reg_entrada[15] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1646 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][17] ) 
    , .D ( sos2_reg_entrada[17] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][17] ) 
    , .D ( sos2_reg_entrada[17] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][17] ) 
    , .D ( sos2_reg_entrada[17] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][17] ) 
    , .D ( sos2_reg_entrada[17] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1648 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][17] ) , .D ( partial_1[17] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1652 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][16] ) 
    , .D ( sos2_reg_entrada[16] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1658 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][16] ) 
    , .D ( sos2_reg_entrada[16] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1646 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][16] ) 
    , .D ( sos2_reg_entrada[16] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[2][18] ) 
    , .D ( sos2_reg_entrada[18] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[1][18] ) 
    , .D ( sos2_reg_entrada[18] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_0_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[0][18] ) 
    , .D ( sos2_reg_entrada[18] ) ) ;
DFFARX1 sos1_reg_pila_registro_reg_7_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1648 ) 
    , .Q ( \sos1_reg/bank_registro_registros[7][18] ) , .D ( partial_1[18] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][17] ) 
    , .D ( sos2_reg_entrada[17] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][17] ) 
    , .D ( sos2_reg_entrada[17] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1652 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][17] ) 
    , .D ( sos2_reg_entrada[17] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1660 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][17] ) 
    , .D ( sos2_reg_entrada[17] ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1648 ) , .QN ( n696 ) 
    , .D ( bajo_reg_entrada[1] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_0_ (.SETB ( n1650 ) 
    , .QN ( bank_registro_registros[16] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n698 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1648 ) , .QN ( n698 ) 
    , .D ( bajo_reg_entrada[0] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[7][18] ) 
    , .D ( sos2_reg_entrada[18] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[6][18] ) 
    , .D ( sos2_reg_entrada[18] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[5][18] ) 
    , .D ( sos2_reg_entrada[18] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[4][18] ) 
    , .D ( sos2_reg_entrada[18] ) ) ;
DFFARX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1648 ) 
    , .Q ( \sos2_reg/bank_registro_registros[3][18] ) 
    , .D ( sos2_reg_entrada[18] ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1646 ) , .QN ( n688 ) 
    , .D ( bajo_reg_entrada[5] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_4_ (.SETB ( n1649 ) 
    , .QN ( bank_registro_registros[20] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n690 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1646 ) , .QN ( n690 ) 
    , .D ( bajo_reg_entrada[4] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_3_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[19] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n692 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1646 ) , .QN ( n692 ) 
    , .D ( bajo_reg_entrada[3] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_2_ (.SETB ( n1650 ) 
    , .QN ( bank_registro_registros[18] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n694 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1648 ) , .QN ( n694 ) 
    , .D ( bajo_reg_entrada[2] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_1_ (.SETB ( n1649 ) 
    , .QN ( bank_registro_registros[17] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n696 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1646 ) , .QN ( n680 ) 
    , .D ( bajo_reg_entrada[9] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_8_ (.SETB ( n1652 ) 
    , .QN ( bank_registro_registros[24] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n682 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1646 ) , .QN ( n682 ) 
    , .D ( bajo_reg_entrada[8] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_7_ (.SETB ( n1651 ) 
    , .QN ( bank_registro_registros[23] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n684 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1646 ) , .QN ( n684 ) 
    , .D ( bajo_reg_entrada[7] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_6_ (.SETB ( n1646 ) 
    , .QN ( bank_registro_registros[22] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n686 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1646 ) , .QN ( n686 ) 
    , .D ( bajo_reg_entrada[6] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_5_ (.SETB ( n1658 ) 
    , .QN ( bank_registro_registros[21] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n688 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1646 ) , .QN ( n672 ) 
    , .D ( bajo_reg_entrada[13] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_12_ (.SETB ( n1661 ) 
    , .QN ( bank_registro_registros[28] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n674 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1646 ) , .QN ( n674 ) 
    , .D ( bajo_reg_entrada[12] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_11_ (.SETB ( n1652 ) 
    , .QN ( bank_registro_registros[27] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n676 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1646 ) , .QN ( n676 ) 
    , .D ( bajo_reg_entrada[11] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_10_ (.SETB ( n1651 ) 
    , .QN ( bank_registro_registros[26] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n678 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1646 ) , .QN ( n678 ) 
    , .D ( bajo_reg_entrada[10] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_9_ (.SETB ( n1662 ) 
    , .QN ( bank_registro_registros[25] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n680 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1655 ) , .QN ( n664 ) 
    , .D ( bajo_reg_entrada[18] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_16_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[32] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n666 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1654 ) , .QN ( n666 ) 
    , .D ( bajo_reg_entrada[16] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_15_ (.SETB ( n1652 ) 
    , .QN ( bank_registro_registros[31] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n668 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1654 ) , .QN ( n668 ) 
    , .D ( bajo_reg_entrada[15] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_14_ (.SETB ( n1653 ) 
    , .QN ( bank_registro_registros[30] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n670 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_0_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia_delay[0] ) , .RSTB ( n1648 ) , .QN ( n670 ) 
    , .D ( bajo_reg_entrada[14] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_13_ (.SETB ( n1651 ) 
    , .QN ( bank_registro_registros[29] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n672 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1654 ) , .QN ( n654 ) 
    , .D ( bajo_reg_entrada[3] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_2_ (.SETB ( n1651 ) 
    , .QN ( bank_registro_registros[36] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n656 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1657 ) , .QN ( n656 ) 
    , .D ( bajo_reg_entrada[2] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_1_ (.SETB ( n1650 ) 
    , .QN ( bank_registro_registros[35] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n658 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1655 ) , .QN ( n658 ) 
    , .D ( bajo_reg_entrada[1] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_0_ (.SETB ( n1652 ) 
    , .QN ( bank_registro_registros[34] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n660 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1655 ) , .QN ( n660 ) 
    , .D ( bajo_reg_entrada[0] ) ) ;
DFFASX1 in_reg_pila_registro_reg_1_registro_tmp_reg_18_ (.SETB ( n1650 ) 
    , .QN ( bank_registro_registros[33] ) , .CLK ( reloj_secuencia[1] ) 
    , .D ( n664 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1656 ) , .QN ( n646 ) 
    , .D ( bajo_reg_entrada[7] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_6_ (.SETB ( n1649 ) 
    , .QN ( bank_registro_registros[40] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n648 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1654 ) , .QN ( n648 ) 
    , .D ( bajo_reg_entrada[6] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_5_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[39] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n650 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1656 ) , .QN ( n650 ) 
    , .D ( bajo_reg_entrada[5] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_4_ (.SETB ( n1658 ) 
    , .QN ( bank_registro_registros[38] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n652 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1654 ) , .QN ( n652 ) 
    , .D ( bajo_reg_entrada[4] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_3_ (.SETB ( n1652 ) 
    , .QN ( bank_registro_registros[37] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n654 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1655 ) , .QN ( n638 ) 
    , .D ( bajo_reg_entrada[11] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_10_ (.SETB ( n1660 ) 
    , .QN ( bank_registro_registros[44] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n640 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1656 ) , .QN ( n640 ) 
    , .D ( bajo_reg_entrada[10] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_9_ (.SETB ( n1646 ) 
    , .QN ( bank_registro_registros[43] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n642 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1656 ) , .QN ( n642 ) 
    , .D ( bajo_reg_entrada[9] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_8_ (.SETB ( n1662 ) 
    , .QN ( bank_registro_registros[42] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n644 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1657 ) , .QN ( n644 ) 
    , .D ( bajo_reg_entrada[8] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_7_ (.SETB ( n1650 ) 
    , .QN ( bank_registro_registros[41] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n646 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1656 ) , .QN ( n630 ) 
    , .D ( bajo_reg_entrada[15] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_14_ (.SETB ( n1652 ) 
    , .QN ( bank_registro_registros[48] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n632 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1657 ) , .QN ( n632 ) 
    , .D ( bajo_reg_entrada[14] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_13_ (.SETB ( n1659 ) 
    , .QN ( bank_registro_registros[47] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n634 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1656 ) , .QN ( n634 ) 
    , .D ( bajo_reg_entrada[13] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_12_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[46] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n636 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1657 ) , .QN ( n636 ) 
    , .D ( bajo_reg_entrada[12] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_11_ (.SETB ( n1652 ) 
    , .QN ( bank_registro_registros[45] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n638 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1654 ) , .QN ( n620 ) 
    , .D ( bajo_reg_entrada[1] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_0_ (.SETB ( n1650 ) 
    , .QN ( bank_registro_registros[52] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n622 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1654 ) , .QN ( n622 ) 
    , .D ( bajo_reg_entrada[0] ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1655 ) , .QN ( n624 ) 
    , .D ( bajo_reg_entrada[18] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_17_ (.SETB ( n1646 ) 
    , .QN ( bank_registro_registros[51] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n624 ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_16_ (.SETB ( n1651 ) 
    , .QN ( bank_registro_registros[50] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n628 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_1_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia_delay[1] ) , .RSTB ( n1654 ) , .QN ( n628 ) 
    , .D ( bajo_reg_entrada[16] ) ) ;
DFFASX1 in_reg_pila_registro_reg_2_registro_tmp_reg_15_ (.SETB ( n1653 ) 
    , .QN ( bank_registro_registros[49] ) , .CLK ( reloj_secuencia[2] ) 
    , .D ( n630 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1656 ) , .QN ( n612 ) 
    , .D ( bajo_reg_entrada[5] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_4_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[56] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n614 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1656 ) , .QN ( n614 ) 
    , .D ( bajo_reg_entrada[4] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_3_ (.SETB ( n1653 ) 
    , .QN ( bank_registro_registros[55] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n616 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1654 ) , .QN ( n616 ) 
    , .D ( bajo_reg_entrada[3] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_2_ (.SETB ( n1649 ) 
    , .QN ( bank_registro_registros[54] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n618 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1656 ) , .QN ( n618 ) 
    , .D ( bajo_reg_entrada[2] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_1_ (.SETB ( n1655 ) 
    , .QN ( bank_registro_registros[53] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n620 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1657 ) , .QN ( n604 ) 
    , .D ( bajo_reg_entrada[9] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_8_ (.SETB ( n1649 ) 
    , .QN ( bank_registro_registros[60] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n606 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1655 ) , .QN ( n606 ) 
    , .D ( bajo_reg_entrada[8] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_7_ (.SETB ( n1650 ) 
    , .QN ( bank_registro_registros[59] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n608 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1657 ) , .QN ( n608 ) 
    , .D ( bajo_reg_entrada[7] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_6_ (.SETB ( n1650 ) 
    , .QN ( bank_registro_registros[58] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n610 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1654 ) , .QN ( n610 ) 
    , .D ( bajo_reg_entrada[6] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_5_ (.SETB ( n1646 ) 
    , .QN ( bank_registro_registros[57] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n612 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1655 ) , .QN ( n596 ) 
    , .D ( bajo_reg_entrada[13] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_12_ (.SETB ( n1646 ) 
    , .QN ( bank_registro_registros[64] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n598 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1654 ) , .QN ( n598 ) 
    , .D ( bajo_reg_entrada[12] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_11_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[63] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n600 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1656 ) , .QN ( n600 ) 
    , .D ( bajo_reg_entrada[11] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_10_ (.SETB ( n1651 ) 
    , .QN ( bank_registro_registros[62] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n602 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1655 ) , .QN ( n602 ) 
    , .D ( bajo_reg_entrada[10] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_9_ (.SETB ( n1653 ) 
    , .QN ( bank_registro_registros[61] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n604 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1657 ) , .QN ( n588 ) 
    , .D ( bajo_reg_entrada[18] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_16_ (.SETB ( n1649 ) 
    , .QN ( bank_registro_registros[68] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n590 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1655 ) , .QN ( n590 ) 
    , .D ( bajo_reg_entrada[16] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_15_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[67] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n592 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1655 ) , .QN ( n592 ) 
    , .D ( bajo_reg_entrada[15] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_14_ (.SETB ( n1650 ) 
    , .QN ( bank_registro_registros[66] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n594 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_2_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia_delay[2] ) , .RSTB ( n1654 ) , .QN ( n594 ) 
    , .D ( bajo_reg_entrada[14] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_13_ (.SETB ( n1651 ) 
    , .QN ( bank_registro_registros[65] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n596 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1653 ) , .QN ( n578 ) 
    , .D ( bajo_reg_entrada[3] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_2_ (.SETB ( n1646 ) 
    , .QN ( bank_registro_registros[72] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n580 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1653 ) , .QN ( n580 ) 
    , .D ( bajo_reg_entrada[2] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_1_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[71] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n582 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1653 ) , .QN ( n582 ) 
    , .D ( bajo_reg_entrada[1] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_0_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[70] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n584 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1656 ) , .QN ( n584 ) 
    , .D ( bajo_reg_entrada[0] ) ) ;
DFFASX1 in_reg_pila_registro_reg_3_registro_tmp_reg_18_ (.SETB ( n1651 ) 
    , .QN ( bank_registro_registros[69] ) , .CLK ( reloj_secuencia[3] ) 
    , .D ( n588 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1653 ) , .QN ( n570 ) 
    , .D ( bajo_reg_entrada[7] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_6_ (.SETB ( n1653 ) 
    , .QN ( bank_registro_registros[76] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n572 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1653 ) , .QN ( n572 ) 
    , .D ( bajo_reg_entrada[6] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_5_ (.SETB ( n1649 ) 
    , .QN ( bank_registro_registros[75] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n574 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1653 ) , .QN ( n574 ) 
    , .D ( bajo_reg_entrada[5] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_4_ (.SETB ( n1663 ) 
    , .QN ( bank_registro_registros[74] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n576 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1653 ) , .QN ( n576 ) 
    , .D ( bajo_reg_entrada[4] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_3_ (.SETB ( n1650 ) 
    , .QN ( bank_registro_registros[73] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n578 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1653 ) , .QN ( n562 ) 
    , .D ( bajo_reg_entrada[11] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_10_ (.SETB ( n1652 ) 
    , .QN ( bank_registro_registros[80] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n564 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1653 ) , .QN ( n564 ) 
    , .D ( bajo_reg_entrada[10] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_9_ (.SETB ( n1650 ) 
    , .QN ( bank_registro_registros[79] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n566 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1653 ) , .QN ( n566 ) 
    , .D ( bajo_reg_entrada[9] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_8_ (.SETB ( n1646 ) 
    , .QN ( bank_registro_registros[78] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n568 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1653 ) , .QN ( n568 ) 
    , .D ( bajo_reg_entrada[8] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_7_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[77] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n570 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1652 ) , .QN ( n554 ) 
    , .D ( bajo_reg_entrada[15] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_14_ (.SETB ( n1646 ) 
    , .QN ( bank_registro_registros[84] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n556 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1652 ) , .QN ( n556 ) 
    , .D ( bajo_reg_entrada[14] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_13_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[83] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n558 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1652 ) , .QN ( n558 ) 
    , .D ( bajo_reg_entrada[13] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_12_ (.SETB ( n1653 ) 
    , .QN ( bank_registro_registros[82] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n560 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1653 ) , .QN ( n560 ) 
    , .D ( bajo_reg_entrada[12] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_11_ (.SETB ( n1649 ) 
    , .QN ( bank_registro_registros[81] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n562 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1652 ) , .QN ( n544 ) 
    , .D ( bajo_reg_entrada[1] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_0_ (.SETB ( n1653 ) 
    , .QN ( bank_registro_registros[88] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n546 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1652 ) , .QN ( n546 ) 
    , .D ( bajo_reg_entrada[0] ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1652 ) , .QN ( n548 ) 
    , .D ( bajo_reg_entrada[18] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_17_ (.SETB ( n1652 ) 
    , .QN ( bank_registro_registros[87] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n548 ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_16_ (.SETB ( n1650 ) 
    , .QN ( bank_registro_registros[86] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n552 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_3_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia_delay[3] ) , .RSTB ( n1652 ) , .QN ( n552 ) 
    , .D ( bajo_reg_entrada[16] ) ) ;
DFFASX1 in_reg_pila_registro_reg_4_registro_tmp_reg_15_ (.SETB ( n1663 ) 
    , .QN ( bank_registro_registros[85] ) , .CLK ( reloj_secuencia[4] ) 
    , .D ( n554 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1651 ) , .QN ( n536 ) 
    , .D ( bajo_reg_entrada[5] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_4_ (.SETB ( n1660 ) 
    , .QN ( bank_registro_registros[92] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n538 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1652 ) , .QN ( n538 ) 
    , .D ( bajo_reg_entrada[4] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_3_ (.SETB ( n1662 ) 
    , .QN ( bank_registro_registros[91] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n540 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1652 ) , .QN ( n540 ) 
    , .D ( bajo_reg_entrada[3] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_2_ (.SETB ( n1646 ) 
    , .QN ( bank_registro_registros[90] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n542 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1652 ) , .QN ( n542 ) 
    , .D ( bajo_reg_entrada[2] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_1_ (.SETB ( n1651 ) 
    , .QN ( bank_registro_registros[89] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n544 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1651 ) , .QN ( n528 ) 
    , .D ( bajo_reg_entrada[9] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_8_ (.SETB ( n1652 ) 
    , .QN ( bank_registro_registros[96] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n530 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1651 ) , .QN ( n530 ) 
    , .D ( bajo_reg_entrada[8] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_7_ (.SETB ( n1651 ) 
    , .QN ( bank_registro_registros[95] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n532 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1651 ) , .QN ( n532 ) 
    , .D ( bajo_reg_entrada[7] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_6_ (.SETB ( n1653 ) 
    , .QN ( bank_registro_registros[94] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n534 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1651 ) , .QN ( n534 ) 
    , .D ( bajo_reg_entrada[6] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_5_ (.SETB ( n1652 ) 
    , .QN ( bank_registro_registros[93] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n536 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1651 ) , .QN ( n520 ) 
    , .D ( bajo_reg_entrada[13] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_12_ (.SETB ( n1646 ) 
    , .QN ( bank_registro_registros[100] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n522 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1651 ) , .QN ( n522 ) 
    , .D ( bajo_reg_entrada[12] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_11_ (.SETB ( n1660 ) 
    , .QN ( bank_registro_registros[99] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n524 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1651 ) , .QN ( n524 ) 
    , .D ( bajo_reg_entrada[11] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_10_ (.SETB ( n1650 ) 
    , .QN ( bank_registro_registros[98] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n526 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1651 ) , .QN ( n526 ) 
    , .D ( bajo_reg_entrada[10] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_9_ (.SETB ( n1649 ) 
    , .QN ( bank_registro_registros[97] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n528 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1661 ) , .QN ( n512 ) 
    , .D ( bajo_reg_entrada[18] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_16_ (.SETB ( n1651 ) 
    , .QN ( bank_registro_registros[104] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n514 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1651 ) , .QN ( n514 ) 
    , .D ( bajo_reg_entrada[16] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_15_ (.SETB ( n1646 ) 
    , .QN ( bank_registro_registros[103] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n516 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1651 ) , .QN ( n516 ) 
    , .D ( bajo_reg_entrada[15] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_14_ (.SETB ( n1649 ) 
    , .QN ( bank_registro_registros[102] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n518 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_4_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia_delay[4] ) , .RSTB ( n1651 ) , .QN ( n518 ) 
    , .D ( bajo_reg_entrada[14] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_13_ (.SETB ( n1652 ) 
    , .QN ( bank_registro_registros[101] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n520 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1653 ) , .QN ( n502 ) 
    , .D ( bajo_reg_entrada[3] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_2_ (.SETB ( n1650 ) 
    , .QN ( bank_registro_registros[108] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n504 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1649 ) , .QN ( n504 ) 
    , .D ( bajo_reg_entrada[2] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_1_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[107] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n506 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1659 ) , .QN ( n506 ) 
    , .D ( bajo_reg_entrada[1] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_0_ (.SETB ( n1661 ) 
    , .QN ( bank_registro_registros[106] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n508 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1662 ) , .QN ( n508 ) 
    , .D ( bajo_reg_entrada[0] ) ) ;
DFFASX1 in_reg_pila_registro_reg_5_registro_tmp_reg_18_ (.SETB ( n1653 ) 
    , .QN ( bank_registro_registros[105] ) , .CLK ( reloj_secuencia[5] ) 
    , .D ( n512 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1652 ) , .QN ( n494 ) 
    , .D ( bajo_reg_entrada[7] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_6_ (.SETB ( n1660 ) 
    , .QN ( bank_registro_registros[112] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n496 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1663 ) , .QN ( n496 ) 
    , .D ( bajo_reg_entrada[6] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_5_ (.SETB ( n1650 ) 
    , .QN ( bank_registro_registros[111] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n498 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1651 ) , .QN ( n498 ) 
    , .D ( bajo_reg_entrada[5] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_4_ (.SETB ( n1649 ) 
    , .QN ( bank_registro_registros[110] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n500 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1646 ) , .QN ( n500 ) 
    , .D ( bajo_reg_entrada[4] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_3_ (.SETB ( n1652 ) 
    , .QN ( bank_registro_registros[109] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n502 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1650 ) , .QN ( n486 ) 
    , .D ( bajo_reg_entrada[11] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_10_ (.SETB ( n1662 ) 
    , .QN ( bank_registro_registros[116] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n488 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1650 ) , .QN ( n488 ) 
    , .D ( bajo_reg_entrada[10] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_9_ (.SETB ( n1663 ) 
    , .QN ( bank_registro_registros[115] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n490 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1647 ) , .QN ( n490 ) 
    , .D ( bajo_reg_entrada[9] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_8_ (.SETB ( n1659 ) 
    , .QN ( bank_registro_registros[114] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n492 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1650 ) , .QN ( n492 ) 
    , .D ( bajo_reg_entrada[8] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_7_ (.SETB ( n1652 ) 
    , .QN ( bank_registro_registros[113] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n494 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1650 ) , .QN ( n478 ) 
    , .D ( bajo_reg_entrada[15] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_14_ (.SETB ( n1663 ) 
    , .QN ( bank_registro_registros[120] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n480 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1650 ) , .QN ( n480 ) 
    , .D ( bajo_reg_entrada[14] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_13_ (.SETB ( n1646 ) 
    , .QN ( bank_registro_registros[119] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n482 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1650 ) , .QN ( n482 ) 
    , .D ( bajo_reg_entrada[13] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_12_ (.SETB ( n1660 ) 
    , .QN ( bank_registro_registros[118] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n484 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1650 ) , .QN ( n484 ) 
    , .D ( bajo_reg_entrada[12] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_11_ (.SETB ( n1661 ) 
    , .QN ( bank_registro_registros[117] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n486 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1650 ) , .QN ( n468 ) 
    , .D ( bajo_reg_entrada[1] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_0_ (.SETB ( n1646 ) 
    , .QN ( bank_registro_registros[124] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n470 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1650 ) , .QN ( n470 ) 
    , .D ( bajo_reg_entrada[0] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_18_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[123] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n472 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1650 ) , .QN ( n472 ) 
    , .D ( bajo_reg_entrada[18] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_16_ (.SETB ( n1662 ) 
    , .QN ( bank_registro_registros[122] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n476 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_5_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia_delay[5] ) , .RSTB ( n1650 ) , .QN ( n476 ) 
    , .D ( bajo_reg_entrada[16] ) ) ;
DFFASX1 in_reg_pila_registro_reg_6_registro_tmp_reg_15_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[121] ) , .CLK ( reloj_secuencia[6] ) 
    , .D ( n478 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1649 ) , .QN ( n460 ) 
    , .D ( bajo_reg_entrada[5] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_4_ (.SETB ( n1661 ) 
    , .QN ( bank_registro_registros[128] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n462 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1649 ) , .QN ( n462 ) 
    , .D ( bajo_reg_entrada[4] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_3_ (.SETB ( n1660 ) 
    , .QN ( bank_registro_registros[127] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n464 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1649 ) , .QN ( n464 ) 
    , .D ( bajo_reg_entrada[3] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_2_ (.SETB ( n1662 ) 
    , .QN ( bank_registro_registros[126] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n466 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1650 ) , .QN ( n466 ) 
    , .D ( bajo_reg_entrada[2] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_1_ (.SETB ( n1659 ) 
    , .QN ( bank_registro_registros[125] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n468 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1649 ) , .QN ( n452 ) 
    , .D ( bajo_reg_entrada[9] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_8_ (.SETB ( n1651 ) 
    , .QN ( bank_registro_registros[132] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n454 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1649 ) , .QN ( n454 ) 
    , .D ( bajo_reg_entrada[8] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_7_ (.SETB ( n1651 ) 
    , .QN ( bank_registro_registros[131] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n456 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1649 ) , .QN ( n456 ) 
    , .D ( bajo_reg_entrada[7] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_6_ (.SETB ( n1646 ) 
    , .QN ( bank_registro_registros[130] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n458 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1649 ) , .QN ( n458 ) 
    , .D ( bajo_reg_entrada[6] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_5_ (.SETB ( n1658 ) 
    , .QN ( bank_registro_registros[129] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n460 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1650 ) , .QN ( n444 ) 
    , .D ( bajo_reg_entrada[13] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_12_ (.SETB ( n1652 ) 
    , .QN ( bank_registro_registros[136] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n446 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1657 ) , .QN ( n446 ) 
    , .D ( bajo_reg_entrada[12] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_11_ (.SETB ( n1653 ) 
    , .QN ( bank_registro_registros[135] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n448 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1652 ) , .QN ( n448 ) 
    , .D ( bajo_reg_entrada[11] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_10_ (.SETB ( n1651 ) 
    , .QN ( bank_registro_registros[134] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n450 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1649 ) , .QN ( n450 ) 
    , .D ( bajo_reg_entrada[10] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_9_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[133] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n452 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1646 ) , .QN ( n436 ) 
    , .D ( bajo_reg_entrada[18] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_16_ (.SETB ( n1658 ) 
    , .QN ( bank_registro_registros[140] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n438 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1649 ) , .QN ( n438 ) 
    , .D ( bajo_reg_entrada[16] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_15_ (.SETB ( n1649 ) 
    , .QN ( bank_registro_registros[139] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n440 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1646 ) , .QN ( n440 ) 
    , .D ( bajo_reg_entrada[15] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_14_ (.SETB ( n1647 ) 
    , .QN ( bank_registro_registros[138] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n442 ) ) ;
DFFARX1 bajo_reg_pila_registro_reg_6_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia_delay[6] ) , .RSTB ( n1647 ) , .QN ( n442 ) 
    , .D ( bajo_reg_entrada[14] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_13_ (.SETB ( n1653 ) 
    , .QN ( bank_registro_registros[137] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n444 ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1653 ) 
    , .Q ( filtro_pipelining_salida[6] ) , .D ( alto_reg_entrada[6] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1661 ) 
    , .Q ( filtro_pipelining_salida[5] ) , .D ( alto_reg_entrada[5] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1658 ) 
    , .Q ( filtro_pipelining_salida[4] ) , .D ( alto_reg_entrada[4] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1652 ) 
    , .Q ( filtro_pipelining_salida[3] ) , .D ( alto_reg_entrada[3] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1649 ) 
    , .Q ( filtro_pipelining_salida[2] ) , .D ( alto_reg_entrada[2] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1660 ) 
    , .Q ( filtro_pipelining_salida[1] ) , .D ( alto_reg_entrada[1] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1659 ) 
    , .Q ( filtro_pipelining_salida[0] ) , .D ( alto_reg_entrada[0] ) ) ;
DFFASX1 in_reg_pila_registro_reg_7_registro_tmp_reg_18_ (.SETB ( n1659 ) 
    , .QN ( bank_registro_registros[141] ) , .CLK ( reloj_secuencia[7] ) 
    , .D ( n436 ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1650 ) 
    , .Q ( filtro_pipelining_salida[14] ) , .D ( alto_reg_entrada[14] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1661 ) 
    , .Q ( filtro_pipelining_salida[13] ) , .D ( alto_reg_entrada[13] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1646 ) 
    , .Q ( filtro_pipelining_salida[12] ) , .D ( alto_reg_entrada[12] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1658 ) 
    , .Q ( filtro_pipelining_salida[11] ) , .D ( alto_reg_entrada[11] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1649 ) 
    , .Q ( filtro_pipelining_salida[10] ) , .D ( alto_reg_entrada[10] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1649 ) 
    , .Q ( filtro_pipelining_salida[9] ) , .D ( alto_reg_entrada[9] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1647 ) 
    , .Q ( filtro_pipelining_salida[8] ) , .D ( alto_reg_entrada[8] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1649 ) 
    , .Q ( filtro_pipelining_salida[7] ) , .D ( alto_reg_entrada[7] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1662 ) 
    , .Q ( filtro_pipelining_salida[22] ) , .D ( alto_reg_entrada[6] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1649 ) 
    , .Q ( filtro_pipelining_salida[21] ) , .D ( alto_reg_entrada[5] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1652 ) 
    , .Q ( filtro_pipelining_salida[20] ) , .D ( alto_reg_entrada[4] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1661 ) 
    , .Q ( filtro_pipelining_salida[19] ) , .D ( alto_reg_entrada[3] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1646 ) 
    , .Q ( filtro_pipelining_salida[18] ) , .D ( alto_reg_entrada[2] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1652 ) 
    , .Q ( filtro_pipelining_salida[17] ) , .D ( alto_reg_entrada[1] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1649 ) 
    , .Q ( filtro_pipelining_salida[16] ) , .D ( alto_reg_entrada[0] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_0_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1646 ) 
    , .Q ( filtro_pipelining_salida[15] ) , .D ( alto_reg_entrada[15] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1652 ) 
    , .Q ( filtro_pipelining_salida[30] ) , .D ( alto_reg_entrada[14] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1662 ) 
    , .Q ( filtro_pipelining_salida[29] ) , .D ( alto_reg_entrada[13] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1647 ) 
    , .Q ( filtro_pipelining_salida[28] ) , .D ( alto_reg_entrada[12] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1658 ) 
    , .Q ( filtro_pipelining_salida[27] ) , .D ( alto_reg_entrada[11] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1652 ) 
    , .Q ( filtro_pipelining_salida[26] ) , .D ( alto_reg_entrada[10] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[25] ) , .D ( alto_reg_entrada[9] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1663 ) 
    , .Q ( filtro_pipelining_salida[24] ) , .D ( alto_reg_entrada[8] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1662 ) 
    , .Q ( filtro_pipelining_salida[23] ) , .D ( alto_reg_entrada[7] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1653 ) 
    , .Q ( filtro_pipelining_salida[38] ) , .D ( alto_reg_entrada[6] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1652 ) 
    , .Q ( filtro_pipelining_salida[37] ) , .D ( alto_reg_entrada[5] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1652 ) 
    , .Q ( filtro_pipelining_salida[36] ) , .D ( alto_reg_entrada[4] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1653 ) 
    , .Q ( filtro_pipelining_salida[35] ) , .D ( alto_reg_entrada[3] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1660 ) 
    , .Q ( filtro_pipelining_salida[34] ) , .D ( alto_reg_entrada[2] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1659 ) 
    , .Q ( filtro_pipelining_salida[33] ) , .D ( alto_reg_entrada[1] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1649 ) 
    , .Q ( filtro_pipelining_salida[32] ) , .D ( alto_reg_entrada[0] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_1_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1653 ) 
    , .Q ( filtro_pipelining_salida[31] ) , .D ( alto_reg_entrada[15] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1647 ) 
    , .Q ( filtro_pipelining_salida[46] ) , .D ( alto_reg_entrada[14] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1646 ) 
    , .Q ( filtro_pipelining_salida[45] ) , .D ( alto_reg_entrada[13] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1658 ) 
    , .Q ( filtro_pipelining_salida[44] ) , .D ( alto_reg_entrada[12] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1653 ) 
    , .Q ( filtro_pipelining_salida[43] ) , .D ( alto_reg_entrada[11] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1646 ) 
    , .Q ( filtro_pipelining_salida[42] ) , .D ( alto_reg_entrada[10] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[41] ) , .D ( alto_reg_entrada[9] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1650 ) 
    , .Q ( filtro_pipelining_salida[40] ) , .D ( alto_reg_entrada[8] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1647 ) 
    , .Q ( filtro_pipelining_salida[39] ) , .D ( alto_reg_entrada[7] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[54] ) , .D ( alto_reg_entrada[6] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1658 ) 
    , .Q ( filtro_pipelining_salida[53] ) , .D ( alto_reg_entrada[5] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1646 ) 
    , .Q ( filtro_pipelining_salida[52] ) , .D ( alto_reg_entrada[4] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1647 ) 
    , .Q ( filtro_pipelining_salida[51] ) , .D ( alto_reg_entrada[3] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[50] ) , .D ( alto_reg_entrada[2] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1650 ) 
    , .Q ( filtro_pipelining_salida[49] ) , .D ( alto_reg_entrada[1] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1659 ) 
    , .Q ( filtro_pipelining_salida[48] ) , .D ( alto_reg_entrada[0] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_2_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[47] ) , .D ( alto_reg_entrada[15] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1647 ) 
    , .Q ( filtro_pipelining_salida[62] ) , .D ( alto_reg_entrada[14] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1646 ) 
    , .Q ( filtro_pipelining_salida[61] ) , .D ( alto_reg_entrada[13] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1646 ) 
    , .Q ( filtro_pipelining_salida[60] ) , .D ( alto_reg_entrada[12] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1646 ) 
    , .Q ( filtro_pipelining_salida[59] ) , .D ( alto_reg_entrada[11] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[58] ) , .D ( alto_reg_entrada[10] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1660 ) 
    , .Q ( filtro_pipelining_salida[57] ) , .D ( alto_reg_entrada[9] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1663 ) 
    , .Q ( filtro_pipelining_salida[56] ) , .D ( alto_reg_entrada[8] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1650 ) 
    , .Q ( filtro_pipelining_salida[55] ) , .D ( alto_reg_entrada[7] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1653 ) 
    , .Q ( filtro_pipelining_salida[70] ) , .D ( alto_reg_entrada[6] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1647 ) 
    , .Q ( filtro_pipelining_salida[69] ) , .D ( alto_reg_entrada[5] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1653 ) 
    , .Q ( filtro_pipelining_salida[68] ) , .D ( alto_reg_entrada[4] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1659 ) 
    , .Q ( filtro_pipelining_salida[67] ) , .D ( alto_reg_entrada[3] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1649 ) 
    , .Q ( filtro_pipelining_salida[66] ) , .D ( alto_reg_entrada[2] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1661 ) 
    , .Q ( filtro_pipelining_salida[65] ) , .D ( alto_reg_entrada[1] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[64] ) , .D ( alto_reg_entrada[0] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_3_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1652 ) 
    , .Q ( filtro_pipelining_salida[63] ) , .D ( alto_reg_entrada[15] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1646 ) 
    , .Q ( filtro_pipelining_salida[78] ) , .D ( alto_reg_entrada[14] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1653 ) 
    , .Q ( filtro_pipelining_salida[77] ) , .D ( alto_reg_entrada[13] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1647 ) 
    , .Q ( filtro_pipelining_salida[76] ) , .D ( alto_reg_entrada[12] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1661 ) 
    , .Q ( filtro_pipelining_salida[75] ) , .D ( alto_reg_entrada[11] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[74] ) , .D ( alto_reg_entrada[10] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[73] ) , .D ( alto_reg_entrada[9] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[72] ) , .D ( alto_reg_entrada[8] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1660 ) 
    , .Q ( filtro_pipelining_salida[71] ) , .D ( alto_reg_entrada[7] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1647 ) 
    , .Q ( filtro_pipelining_salida[86] ) , .D ( alto_reg_entrada[6] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1649 ) 
    , .Q ( filtro_pipelining_salida[85] ) , .D ( alto_reg_entrada[5] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1647 ) 
    , .Q ( filtro_pipelining_salida[84] ) , .D ( alto_reg_entrada[4] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[83] ) , .D ( alto_reg_entrada[3] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1652 ) 
    , .Q ( filtro_pipelining_salida[82] ) , .D ( alto_reg_entrada[2] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1649 ) 
    , .Q ( filtro_pipelining_salida[81] ) , .D ( alto_reg_entrada[1] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1650 ) 
    , .Q ( filtro_pipelining_salida[80] ) , .D ( alto_reg_entrada[0] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_4_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1650 ) 
    , .Q ( filtro_pipelining_salida[79] ) , .D ( alto_reg_entrada[15] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1649 ) 
    , .Q ( filtro_pipelining_salida[94] ) , .D ( alto_reg_entrada[14] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1649 ) 
    , .Q ( filtro_pipelining_salida[93] ) , .D ( alto_reg_entrada[13] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1653 ) 
    , .Q ( filtro_pipelining_salida[92] ) , .D ( alto_reg_entrada[12] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1650 ) 
    , .Q ( filtro_pipelining_salida[91] ) , .D ( alto_reg_entrada[11] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1659 ) 
    , .Q ( filtro_pipelining_salida[90] ) , .D ( alto_reg_entrada[10] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1650 ) 
    , .Q ( filtro_pipelining_salida[89] ) , .D ( alto_reg_entrada[9] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1658 ) 
    , .Q ( filtro_pipelining_salida[88] ) , .D ( alto_reg_entrada[8] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[87] ) , .D ( alto_reg_entrada[7] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1660 ) 
    , .Q ( filtro_pipelining_salida[102] ) , .D ( alto_reg_entrada[6] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1660 ) 
    , .Q ( filtro_pipelining_salida[101] ) , .D ( alto_reg_entrada[5] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1653 ) 
    , .Q ( filtro_pipelining_salida[100] ) , .D ( alto_reg_entrada[4] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[99] ) , .D ( alto_reg_entrada[3] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[98] ) , .D ( alto_reg_entrada[2] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1647 ) 
    , .Q ( filtro_pipelining_salida[97] ) , .D ( alto_reg_entrada[1] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1650 ) 
    , .Q ( filtro_pipelining_salida[96] ) , .D ( alto_reg_entrada[0] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_5_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1652 ) 
    , .Q ( filtro_pipelining_salida[95] ) , .D ( alto_reg_entrada[15] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1653 ) 
    , .Q ( filtro_pipelining_salida[110] ) , .D ( alto_reg_entrada[14] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1662 ) 
    , .Q ( filtro_pipelining_salida[109] ) , .D ( alto_reg_entrada[13] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[108] ) , .D ( alto_reg_entrada[12] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1650 ) 
    , .Q ( filtro_pipelining_salida[107] ) , .D ( alto_reg_entrada[11] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1658 ) 
    , .Q ( filtro_pipelining_salida[106] ) , .D ( alto_reg_entrada[10] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1652 ) 
    , .Q ( filtro_pipelining_salida[105] ) , .D ( alto_reg_entrada[9] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1659 ) 
    , .Q ( filtro_pipelining_salida[104] ) , .D ( alto_reg_entrada[8] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1662 ) 
    , .Q ( filtro_pipelining_salida[103] ) , .D ( alto_reg_entrada[7] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1653 ) 
    , .Q ( filtro_pipelining_salida[118] ) , .D ( alto_reg_entrada[6] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1646 ) 
    , .Q ( filtro_pipelining_salida[117] ) , .D ( alto_reg_entrada[5] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1652 ) 
    , .Q ( filtro_pipelining_salida[116] ) , .D ( alto_reg_entrada[4] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1646 ) 
    , .Q ( filtro_pipelining_salida[115] ) , .D ( alto_reg_entrada[3] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1662 ) 
    , .Q ( filtro_pipelining_salida[114] ) , .D ( alto_reg_entrada[2] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1647 ) 
    , .Q ( filtro_pipelining_salida[113] ) , .D ( alto_reg_entrada[1] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1652 ) 
    , .Q ( filtro_pipelining_salida[112] ) , .D ( alto_reg_entrada[0] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_6_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1661 ) 
    , .Q ( filtro_pipelining_salida[111] ) , .D ( alto_reg_entrada[15] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1663 ) 
    , .Q ( filtro_pipelining_salida[126] ) , .D ( alto_reg_entrada[14] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1663 ) 
    , .Q ( filtro_pipelining_salida[125] ) , .D ( alto_reg_entrada[13] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1661 ) 
    , .Q ( filtro_pipelining_salida[124] ) , .D ( alto_reg_entrada[12] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1662 ) 
    , .Q ( filtro_pipelining_salida[123] ) , .D ( alto_reg_entrada[11] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1661 ) 
    , .Q ( filtro_pipelining_salida[122] ) , .D ( alto_reg_entrada[10] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1649 ) 
    , .Q ( filtro_pipelining_salida[121] ) , .D ( alto_reg_entrada[9] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1659 ) 
    , .Q ( filtro_pipelining_salida[120] ) , .D ( alto_reg_entrada[8] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1649 ) 
    , .Q ( filtro_pipelining_salida[119] ) , .D ( alto_reg_entrada[7] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1649 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][6] ) , .D ( partial_2_L[6] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][5] ) , .D ( partial_2_L[5] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][4] ) , .D ( partial_2_L[4] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][3] ) , .D ( partial_2_L[3] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][2] ) , .D ( partial_2_L[2] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][1] ) , .D ( partial_2_L[1] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][0] ) , .D ( partial_2_L[0] ) ) ;
DFFARX1 alto_reg_pila_registro_reg_7_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1651 ) 
    , .Q ( filtro_pipelining_salida[127] ) , .D ( alto_reg_entrada[15] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][14] ) , .D ( partial_2_L[14] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][13] ) , .D ( partial_2_L[13] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][12] ) , .D ( partial_2_L[12] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][11] ) , .D ( partial_2_L[11] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1646 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][10] ) , .D ( partial_2_L[10] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1652 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][9] ) , .D ( partial_2_L[9] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][8] ) , .D ( partial_2_L[8] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1647 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][7] ) , .D ( partial_2_L[7] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][3] ) , .D ( partial_2_L[3] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][2] ) , .D ( partial_2_L[2] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][1] ) , .D ( partial_2_L[1] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][0] ) , .D ( partial_2_L[0] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1646 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][18] ) , .D ( partial_2_L[18] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][17] ) , .D ( partial_2_L[17] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1646 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][16] ) , .D ( partial_2_L[16] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_0_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1652 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[0][15] ) , .D ( partial_2_L[15] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][11] ) , .D ( partial_2_L[11] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][10] ) , .D ( partial_2_L[10] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][9] ) , .D ( partial_2_L[9] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][8] ) , .D ( partial_2_L[8] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][7] ) , .D ( partial_2_L[7] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][6] ) , .D ( partial_2_L[6] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][5] ) , .D ( partial_2_L[5] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][4] ) , .D ( partial_2_L[4] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][0] ) , .D ( partial_2_L[0] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][18] ) , .D ( partial_2_L[18] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][17] ) , .D ( partial_2_L[17] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][16] ) , .D ( partial_2_L[16] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][15] ) , .D ( partial_2_L[15] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][14] ) , .D ( partial_2_L[14] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][13] ) , .D ( partial_2_L[13] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_1_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[1][12] ) , .D ( partial_2_L[12] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][8] ) , .D ( partial_2_L[8] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][7] ) , .D ( partial_2_L[7] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][6] ) , .D ( partial_2_L[6] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][5] ) , .D ( partial_2_L[5] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][4] ) , .D ( partial_2_L[4] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][3] ) , .D ( partial_2_L[3] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][2] ) , .D ( partial_2_L[2] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][1] ) , .D ( partial_2_L[1] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][16] ) , .D ( partial_2_L[16] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][15] ) , .D ( partial_2_L[15] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][14] ) , .D ( partial_2_L[14] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][13] ) , .D ( partial_2_L[13] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][12] ) , .D ( partial_2_L[12] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][11] ) , .D ( partial_2_L[11] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][10] ) , .D ( partial_2_L[10] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][9] ) , .D ( partial_2_L[9] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][5] ) , .D ( partial_2_L[5] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][4] ) , .D ( partial_2_L[4] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][3] ) , .D ( partial_2_L[3] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][2] ) , .D ( partial_2_L[2] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][1] ) , .D ( partial_2_L[1] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][0] ) , .D ( partial_2_L[0] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][18] ) , .D ( partial_2_L[18] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_2_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[2][17] ) , .D ( partial_2_L[17] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][13] ) , .D ( partial_2_L[13] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][12] ) , .D ( partial_2_L[12] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][11] ) , .D ( partial_2_L[11] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][10] ) , .D ( partial_2_L[10] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][9] ) , .D ( partial_2_L[9] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][8] ) , .D ( partial_2_L[8] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][7] ) , .D ( partial_2_L[7] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][6] ) , .D ( partial_2_L[6] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][2] ) , .D ( partial_2_L[2] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][1] ) , .D ( partial_2_L[1] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][0] ) , .D ( partial_2_L[0] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][18] ) , .D ( partial_2_L[18] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][17] ) , .D ( partial_2_L[17] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][16] ) , .D ( partial_2_L[16] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][15] ) , .D ( partial_2_L[15] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_3_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[3][14] ) , .D ( partial_2_L[14] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][10] ) , .D ( partial_2_L[10] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][9] ) , .D ( partial_2_L[9] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][8] ) , .D ( partial_2_L[8] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][7] ) , .D ( partial_2_L[7] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][6] ) , .D ( partial_2_L[6] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][5] ) , .D ( partial_2_L[5] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][4] ) , .D ( partial_2_L[4] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][3] ) , .D ( partial_2_L[3] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][18] ) , .D ( partial_2_L[18] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][17] ) , .D ( partial_2_L[17] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][16] ) , .D ( partial_2_L[16] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][15] ) , .D ( partial_2_L[15] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][14] ) , .D ( partial_2_L[14] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][13] ) , .D ( partial_2_L[13] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][12] ) , .D ( partial_2_L[12] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_4_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[4][11] ) , .D ( partial_2_L[11] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][7] ) , .D ( partial_2_L[7] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][6] ) , .D ( partial_2_L[6] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][5] ) , .D ( partial_2_L[5] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][4] ) , .D ( partial_2_L[4] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][3] ) , .D ( partial_2_L[3] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][2] ) , .D ( partial_2_L[2] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][1] ) , .D ( partial_2_L[1] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][0] ) , .D ( partial_2_L[0] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][15] ) , .D ( partial_2_L[15] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][14] ) , .D ( partial_2_L[14] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][13] ) , .D ( partial_2_L[13] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][12] ) , .D ( partial_2_L[12] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][11] ) , .D ( partial_2_L[11] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][10] ) , .D ( partial_2_L[10] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][9] ) , .D ( partial_2_L[9] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][8] ) , .D ( partial_2_L[8] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][4] ) , .D ( partial_2_L[4] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][3] ) , .D ( partial_2_L[3] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][2] ) , .D ( partial_2_L[2] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][1] ) , .D ( partial_2_L[1] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][0] ) , .D ( partial_2_L[0] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][18] ) , .D ( partial_2_L[18] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][17] ) , .D ( partial_2_L[17] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_5_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[5][16] ) , .D ( partial_2_L[16] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][12] ) , .D ( partial_2_L[12] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][11] ) , .D ( partial_2_L[11] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][10] ) , .D ( partial_2_L[10] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][9] ) , .D ( partial_2_L[9] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][8] ) , .D ( partial_2_L[8] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][7] ) , .D ( partial_2_L[7] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][6] ) , .D ( partial_2_L[6] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][5] ) , .D ( partial_2_L[5] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][1] ) , .D ( partial_2_L[1] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][0] ) , .D ( partial_2_L[0] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][18] ) , .D ( partial_2_L[18] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][17] ) , .D ( partial_2_L[17] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][16] ) , .D ( partial_2_L[16] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][15] ) , .D ( partial_2_L[15] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][14] ) , .D ( partial_2_L[14] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_6_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[6][13] ) , .D ( partial_2_L[13] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][9] ) , .D ( partial_2_L[9] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][8] ) , .D ( partial_2_L[8] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][7] ) , .D ( partial_2_L[7] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][6] ) , .D ( partial_2_L[6] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][5] ) , .D ( partial_2_L[5] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][4] ) , .D ( partial_2_L[4] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][3] ) , .D ( partial_2_L[3] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][2] ) , .D ( partial_2_L[2] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][17] ) , .D ( partial_2_L[17] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][16] ) , .D ( partial_2_L[16] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][15] ) , .D ( partial_2_L[15] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][14] ) , .D ( partial_2_L[14] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][13] ) , .D ( partial_2_L[13] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][12] ) , .D ( partial_2_L[12] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][11] ) , .D ( partial_2_L[11] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][10] ) , .D ( partial_2_L[10] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][6] ) , .D ( partial_2_H[6] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][5] ) , .D ( partial_2_H[5] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][4] ) , .D ( partial_2_H[4] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][3] ) , .D ( partial_2_H[3] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][2] ) , .D ( partial_2_H[2] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][1] ) , .D ( partial_2_H[1] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][0] ) , .D ( partial_2_H[0] ) ) ;
DFFARX1 pos_L_reg_pila_registro_reg_7_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_L_reg/bank_registro_registros[7][18] ) , .D ( partial_2_L[18] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][14] ) , .D ( partial_2_H[14] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][13] ) , .D ( partial_2_H[13] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][12] ) , .D ( partial_2_H[12] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1652 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][11] ) , .D ( partial_2_H[11] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][10] ) , .D ( partial_2_H[10] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][9] ) , .D ( partial_2_H[9] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][8] ) , .D ( partial_2_H[8] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][7] ) , .D ( partial_2_H[7] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][3] ) , .D ( partial_2_H[3] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1652 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][2] ) , .D ( partial_2_H[2] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1647 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][1] ) , .D ( partial_2_H[1] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][0] ) , .D ( partial_2_H[0] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][18] ) , .D ( partial_2_H[18] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][17] ) , .D ( partial_2_H[17] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][16] ) , .D ( partial_2_H[16] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_0_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[0] ) , .RSTB ( n1646 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[0][15] ) , .D ( partial_2_H[15] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][11] ) , .D ( partial_2_H[11] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1646 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][10] ) , .D ( partial_2_H[10] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][9] ) , .D ( partial_2_H[9] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][8] ) , .D ( partial_2_H[8] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1647 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][7] ) , .D ( partial_2_H[7] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][6] ) , .D ( partial_2_H[6] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][5] ) , .D ( partial_2_H[5] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1652 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][4] ) , .D ( partial_2_H[4] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1651 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][0] ) , .D ( partial_2_H[0] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][18] ) , .D ( partial_2_H[18] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][17] ) , .D ( partial_2_H[17] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1647 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][16] ) , .D ( partial_2_H[16] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1649 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][15] ) , .D ( partial_2_H[15] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1649 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][14] ) , .D ( partial_2_H[14] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1646 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][13] ) , .D ( partial_2_H[13] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_1_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[1] ) , .RSTB ( n1646 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[1][12] ) , .D ( partial_2_H[12] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1651 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][8] ) , .D ( partial_2_H[8] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1649 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][7] ) , .D ( partial_2_H[7] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1646 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][6] ) , .D ( partial_2_H[6] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1647 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][5] ) , .D ( partial_2_H[5] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1651 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][4] ) , .D ( partial_2_H[4] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1647 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][3] ) , .D ( partial_2_H[3] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][2] ) , .D ( partial_2_H[2] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][1] ) , .D ( partial_2_H[1] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][16] ) , .D ( partial_2_H[16] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1651 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][15] ) , .D ( partial_2_H[15] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1652 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][14] ) , .D ( partial_2_H[14] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][13] ) , .D ( partial_2_H[13] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][12] ) , .D ( partial_2_H[12] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][11] ) , .D ( partial_2_H[11] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1647 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][10] ) , .D ( partial_2_H[10] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][9] ) , .D ( partial_2_H[9] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][5] ) , .D ( partial_2_H[5] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1646 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][4] ) , .D ( partial_2_H[4] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1652 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][3] ) , .D ( partial_2_H[3] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][2] ) , .D ( partial_2_H[2] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1646 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][1] ) , .D ( partial_2_H[1] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1652 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][0] ) , .D ( partial_2_H[0] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1651 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][18] ) , .D ( partial_2_H[18] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_2_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[2] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[2][17] ) , .D ( partial_2_H[17] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1649 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][13] ) , .D ( partial_2_H[13] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1651 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][12] ) , .D ( partial_2_H[12] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1649 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][11] ) , .D ( partial_2_H[11] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1646 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][10] ) , .D ( partial_2_H[10] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][9] ) , .D ( partial_2_H[9] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][8] ) , .D ( partial_2_H[8] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][7] ) , .D ( partial_2_H[7] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1649 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][6] ) , .D ( partial_2_H[6] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][2] ) , .D ( partial_2_H[2] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1649 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][1] ) , .D ( partial_2_H[1] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1647 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][0] ) , .D ( partial_2_H[0] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1651 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][18] ) , .D ( partial_2_H[18] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1649 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][17] ) , .D ( partial_2_H[17] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][16] ) , .D ( partial_2_H[16] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][15] ) , .D ( partial_2_H[15] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_3_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[3] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[3][14] ) , .D ( partial_2_H[14] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][10] ) , .D ( partial_2_H[10] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][9] ) , .D ( partial_2_H[9] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1652 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][8] ) , .D ( partial_2_H[8] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1647 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][7] ) , .D ( partial_2_H[7] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1651 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][6] ) , .D ( partial_2_H[6] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][5] ) , .D ( partial_2_H[5] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1646 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][4] ) , .D ( partial_2_H[4] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][3] ) , .D ( partial_2_H[3] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1651 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][18] ) , .D ( partial_2_H[18] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][17] ) , .D ( partial_2_H[17] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1652 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][16] ) , .D ( partial_2_H[16] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][15] ) , .D ( partial_2_H[15] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][14] ) , .D ( partial_2_H[14] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][13] ) , .D ( partial_2_H[13] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1647 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][12] ) , .D ( partial_2_H[12] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_4_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[4] ) , .RSTB ( n1652 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[4][11] ) , .D ( partial_2_H[11] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1649 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][7] ) , .D ( partial_2_H[7] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1658 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][6] ) , .D ( partial_2_H[6] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1646 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][5] ) , .D ( partial_2_H[5] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1647 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][4] ) , .D ( partial_2_H[4] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1647 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][3] ) , .D ( partial_2_H[3] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1649 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][2] ) , .D ( partial_2_H[2] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1646 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][1] ) , .D ( partial_2_H[1] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1649 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][0] ) , .D ( partial_2_H[0] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1651 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][15] ) , .D ( partial_2_H[15] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][14] ) , .D ( partial_2_H[14] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][13] ) , .D ( partial_2_H[13] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1647 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][12] ) , .D ( partial_2_H[12] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1661 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][11] ) , .D ( partial_2_H[11] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1651 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][10] ) , .D ( partial_2_H[10] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1660 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][9] ) , .D ( partial_2_H[9] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][8] ) , .D ( partial_2_H[8] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][4] ) , .D ( partial_2_H[4] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1649 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][3] ) , .D ( partial_2_H[3] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1652 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][2] ) , .D ( partial_2_H[2] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1652 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][1] ) , .D ( partial_2_H[1] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][0] ) , .D ( partial_2_H[0] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1659 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][18] ) , .D ( partial_2_H[18] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1649 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][17] ) , .D ( partial_2_H[17] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_5_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[5] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[5][16] ) , .D ( partial_2_H[16] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1646 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][12] ) , .D ( partial_2_H[12] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1651 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][11] ) , .D ( partial_2_H[11] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][10] ) , .D ( partial_2_H[10] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1652 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][9] ) , .D ( partial_2_H[9] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1647 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][8] ) , .D ( partial_2_H[8] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][7] ) , .D ( partial_2_H[7] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][6] ) , .D ( partial_2_H[6] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1652 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][5] ) , .D ( partial_2_H[5] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_1_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][1] ) , .D ( partial_2_H[1] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_0_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][0] ) , .D ( partial_2_H[0] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][18] ) , .D ( partial_2_H[18] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][17] ) , .D ( partial_2_H[17] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][16] ) , .D ( partial_2_H[16] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][15] ) , .D ( partial_2_H[15] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][14] ) , .D ( partial_2_H[14] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_6_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[6] ) , .RSTB ( n1650 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[6][13] ) , .D ( partial_2_H[13] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_9_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][9] ) , .D ( partial_2_H[9] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_8_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][8] ) , .D ( partial_2_H[8] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_7_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][7] ) , .D ( partial_2_H[7] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_6_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][6] ) , .D ( partial_2_H[6] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_5_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][5] ) , .D ( partial_2_H[5] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_4_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][4] ) , .D ( partial_2_H[4] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_3_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][3] ) , .D ( partial_2_H[3] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_2_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][2] ) , .D ( partial_2_H[2] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_17_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][17] ) , .D ( partial_2_H[17] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_16_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][16] ) , .D ( partial_2_H[16] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_15_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][15] ) , .D ( partial_2_H[15] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_14_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][14] ) , .D ( partial_2_H[14] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_13_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][13] ) , .D ( partial_2_H[13] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_12_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][12] ) , .D ( partial_2_H[12] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_11_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1662 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][11] ) , .D ( partial_2_H[11] ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_10_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1663 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][10] ) , .D ( partial_2_H[10] ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U35 (.A ( n1616 ) , .B ( partial_3_H[18] ) 
    , .CI ( DP_OP_1004J1_67_3033_n53 ) , .CO ( DP_OP_1004J1_67_3033_n45 ) 
    , .S ( DP_OP_1004J1_67_3033_n46 ) ) ;
NAND4X0 U109 (.IN1 ( reloj_secuencia[0] ) , .QN ( n1120 ) 
    , .IN2 ( reloj_secuencia[1] ) , .IN3 ( reloj_secuencia[2] ) 
    , .IN4 ( reloj_secuencia[3] ) ) ;
AND2X1 U108 (.IN1 ( n1033 ) , .IN2 ( reloj_secuencia[4] ) , .Q ( n1125 ) ) ;
NAND2X0 U107 (.IN1 ( reloj_secuencia[0] ) , .IN2 ( reloj_secuencia[1] ) 
    , .QN ( n1121 ) ) ;
AO221X1 U106 (.IN5 ( n1121 ) , .Q ( n1124 ) , .IN2 ( n1034 ) , .IN1 ( n1125 ) 
    , .IN3 ( n1125 ) , .IN4 ( reloj_secuencia[6] ) ) ;
NAND2X0 U105 (.IN1 ( reloj_secuencia[0] ) , .IN2 ( n1124 ) , .QN ( n1122 ) ) ;
NAND4X0 U104 (.IN1 ( reloj_secuencia[1] ) , .QN ( n1123 ) 
    , .IN2 ( reloj_secuencia[2] ) , .IN3 ( reloj_secuencia[0] ) , .IN4 ( n1120 ) ) ;
DFFARX1 pos_H_reg_pila_registro_reg_7_registro_tmp_reg_18_ (
    .CLK ( reloj_secuencia[7] ) , .RSTB ( n1653 ) 
    , .Q ( \pos_H_reg/bank_registro_registros[7][18] ) , .D ( partial_2_H[18] ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U11 (.A ( DP_OP_1004J1_67_3033_n43 ) 
    , .B ( DP_OP_1004J1_67_3033_n40 ) , .CI ( DP_OP_1004J1_67_3033_n11 ) 
    , .CO ( DP_OP_1004J1_67_3033_n10 ) , .S ( alto_reg_entrada[8] ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U12 (.A ( DP_OP_1004J1_67_3033_n49 ) 
    , .B ( DP_OP_1004J1_67_3033_n44 ) , .CI ( DP_OP_1004J1_67_3033_n12 ) 
    , .CO ( DP_OP_1004J1_67_3033_n11 ) , .S ( alto_reg_entrada[7] ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U13 (.A ( DP_OP_1004J1_67_3033_n55 ) 
    , .B ( DP_OP_1004J1_67_3033_n50 ) , .CI ( DP_OP_1004J1_67_3033_n13 ) 
    , .CO ( DP_OP_1004J1_67_3033_n12 ) , .S ( alto_reg_entrada[6] ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U14 (.A ( DP_OP_1004J1_67_3033_n61 ) 
    , .B ( DP_OP_1004J1_67_3033_n56 ) , .CI ( DP_OP_1004J1_67_3033_n14 ) 
    , .CO ( DP_OP_1004J1_67_3033_n13 ) , .S ( alto_reg_entrada[5] ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U40 (.A ( DP_OP_1004J1_67_3033_n60 ) 
    , .B ( DP_OP_1004J1_67_3033_n63 ) , .CI ( DP_OP_1004J1_67_3033_n58 ) 
    , .CO ( DP_OP_1004J1_67_3033_n55 ) , .S ( DP_OP_1004J1_67_3033_n56 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U37 (.A ( DP_OP_1004J1_67_3033_n54 ) 
    , .B ( DP_OP_1004J1_67_3033_n57 ) , .CI ( DP_OP_1004J1_67_3033_n52 ) 
    , .CO ( DP_OP_1004J1_67_3033_n49 ) , .S ( DP_OP_1004J1_67_3033_n50 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U34 (.A ( DP_OP_1004J1_67_3033_n48 ) 
    , .B ( DP_OP_1004J1_67_3033_n51 ) , .CI ( DP_OP_1004J1_67_3033_n46 ) 
    , .CO ( DP_OP_1004J1_67_3033_n43 ) , .S ( DP_OP_1004J1_67_3033_n44 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U32 (.A ( DP_OP_1004J1_67_3033_n47 ) 
    , .B ( DP_OP_1004J1_67_3033_n42 ) , .CI ( DP_OP_1004J1_67_3033_n45 ) 
    , .CO ( DP_OP_1004J1_67_3033_n39 ) , .S ( DP_OP_1004J1_67_3033_n40 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U46 (.A ( DP_OP_1004J1_67_3033_n75 ) 
    , .B ( DP_OP_1004J1_67_3033_n72 ) , .CI ( DP_OP_1004J1_67_3033_n70 ) 
    , .CO ( DP_OP_1004J1_67_3033_n67 ) , .S ( DP_OP_1004J1_67_3033_n68 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U47 (.A ( n1622 ) , .B ( n1614 ) 
    , .CI ( DP_OP_1004J1_67_3033_n77 ) , .CO ( DP_OP_1004J1_67_3033_n69 ) 
    , .S ( DP_OP_1004J1_67_3033_n70 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U39 (.A ( partial_3_H[17] ) 
    , .B ( partial_3_H[8] ) , .CI ( n1619 ) , .CO ( DP_OP_1004J1_67_3033_n53 ) 
    , .S ( DP_OP_1004J1_67_3033_n54 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U15 (.A ( DP_OP_1004J1_67_3033_n67 ) 
    , .B ( DP_OP_1004J1_67_3033_n62 ) , .CI ( DP_OP_1004J1_67_3033_n15 ) 
    , .CO ( DP_OP_1004J1_67_3033_n14 ) , .S ( alto_reg_entrada[4] ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U43 (.A ( DP_OP_1004J1_67_3033_n69 ) 
    , .B ( DP_OP_1004J1_67_3033_n66 ) , .CI ( DP_OP_1004J1_67_3033_n64 ) 
    , .CO ( DP_OP_1004J1_67_3033_n61 ) , .S ( DP_OP_1004J1_67_3033_n62 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U44 (.A ( n1621 ) , .B ( n1613 ) 
    , .CI ( DP_OP_1004J1_67_3033_n71 ) , .CO ( DP_OP_1004J1_67_3033_n63 ) 
    , .S ( DP_OP_1004J1_67_3033_n64 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U36 (.A ( partial_3_H[9] ) , .B ( n1613 ) 
    , .CI ( n1618 ) , .CO ( DP_OP_1004J1_67_3033_n47 ) 
    , .S ( DP_OP_1004J1_67_3033_n48 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U24 (.A ( partial_3_H[15] ) , .B ( n1613 ) 
    , .CI ( partial_3_H[18] ) , .CO ( DP_OP_1004J1_67_3033_n23 ) 
    , .S ( DP_OP_1004J1_67_3033_n24 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U54 (.A ( partial_3_H[3] ) , .B ( n1622 ) 
    , .CI ( n1618 ) , .CO ( DP_OP_1004J1_67_3033_n81 ) 
    , .S ( DP_OP_1004J1_67_3033_n82 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U19 (.A ( n1625 ) , .B ( n1617 ) 
    , .CI ( DP_OP_1004J1_67_3033_n84 ) , .CO ( DP_OP_1004J1_67_3033_n18 ) 
    , .S ( alto_reg_entrada[0] ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U53 (.A ( n1624 ) , .B ( n1616 ) 
    , .CI ( DP_OP_1004J1_67_3033_n83 ) , .CO ( DP_OP_1004J1_67_3033_n79 ) 
    , .S ( DP_OP_1004J1_67_3033_n80 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U49 (.A ( DP_OP_1004J1_67_3033_n81 ) 
    , .B ( DP_OP_1004J1_67_3033_n78 ) , .CI ( DP_OP_1004J1_67_3033_n76 ) 
    , .CO ( DP_OP_1004J1_67_3033_n73 ) , .S ( DP_OP_1004J1_67_3033_n74 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U50 (.A ( n1617 ) , .B ( n1615 ) , .CI ( n1623 ) 
    , .CO ( DP_OP_1004J1_67_3033_n75 ) , .S ( DP_OP_1004J1_67_3033_n76 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U42 (.A ( partial_3_H[16] ) 
    , .B ( partial_3_H[7] ) , .CI ( n1620 ) , .CO ( DP_OP_1004J1_67_3033_n59 ) 
    , .S ( DP_OP_1004J1_67_3033_n60 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U27 (.A ( partial_3_H[13] ) , .B ( n1614 ) 
    , .CI ( n1615 ) , .CO ( DP_OP_1004J1_67_3033_n29 ) 
    , .S ( DP_OP_1004J1_67_3033_n30 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U16 (.A ( DP_OP_1004J1_67_3033_n73 ) 
    , .B ( DP_OP_1004J1_67_3033_n68 ) , .CI ( DP_OP_1004J1_67_3033_n16 ) 
    , .CO ( DP_OP_1004J1_67_3033_n15 ) , .S ( alto_reg_entrada[3] ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U39 (.A ( partial_3_L[15] ) 
    , .B ( partial_3_L[7] ) , .CI ( n1605 ) , .CO ( DP_OP_1003J1_66_5789_n53 ) 
    , .S ( DP_OP_1003J1_66_5789_n54 ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U33 (.A ( partial_3_L[10] ) 
    , .B ( partial_3_L[15] ) , .CI ( n1604 ) , .CO ( DP_OP_1003J1_66_5789_n41 ) 
    , .S ( DP_OP_1003J1_66_5789_n42 ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U37 (.A ( partial_3_L[16] ) 
    , .B ( partial_3_L[8] ) , .CI ( n1604 ) , .CO ( DP_OP_1003J1_66_5789_n49 ) 
    , .S ( DP_OP_1003J1_66_5789_n50 ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U30 (.A ( n1602 ) 
    , .B ( DP_OP_1003J1_66_5789_n41 ) , .CI ( DP_OP_1003J1_66_5789_n38 ) 
    , .CO ( DP_OP_1003J1_66_5789_n35 ) , .S ( DP_OP_1003J1_66_5789_n36 ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U35 (.A ( partial_3_L[17] ) 
    , .B ( partial_3_L[9] ) , .CI ( n1603 ) , .CO ( DP_OP_1003J1_66_5789_n45 ) 
    , .S ( DP_OP_1003J1_66_5789_n46 ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U29 (.A ( partial_3_L[12] ) 
    , .B ( partial_3_L[17] ) , .CI ( n1602 ) , .CO ( DP_OP_1003J1_66_5789_n33 ) 
    , .S ( DP_OP_1003J1_66_5789_n34 ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U32 (.A ( n1599 ) 
    , .B ( DP_OP_1003J1_66_5789_n45 ) , .CI ( DP_OP_1003J1_66_5789_n42 ) 
    , .CO ( DP_OP_1003J1_66_5789_n39 ) , .S ( DP_OP_1003J1_66_5789_n40 ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U55 (.A ( partial_3_H[2] ) , .B ( n1623 ) 
    , .CI ( n1619 ) , .CO ( DP_OP_1004J1_67_3033_n83 ) 
    , .S ( DP_OP_1004J1_67_3033_n84 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U130 (.A ( DP_OP_1002J1_65_247_n186 ) 
    , .B ( DP_OP_1002J1_65_247_n185 ) , .CI ( DP_OP_1002J1_65_247_n165 ) 
    , .CO ( DP_OP_1002J1_65_247_n164 ) , .S ( DP_OP_1002J1_65_247_n272 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U131 (.A ( DP_OP_1002J1_65_247_n188 ) 
    , .B ( DP_OP_1002J1_65_247_n187 ) , .CI ( DP_OP_1002J1_65_247_n166 ) 
    , .CO ( DP_OP_1002J1_65_247_n165 ) , .S ( DP_OP_1002J1_65_247_n271 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U132 (.A ( DP_OP_1002J1_65_247_n190 ) 
    , .B ( DP_OP_1002J1_65_247_n189 ) , .CI ( DP_OP_1002J1_65_247_n167 ) 
    , .CO ( DP_OP_1002J1_65_247_n166 ) , .S ( DP_OP_1002J1_65_247_n270 ) ) ;
HADDX1 DP_OP_1003J1_66_5789_U49 (.B0 ( partial_3_L[10] ) 
    , .A0 ( partial_3_L[2] ) , .C1 ( DP_OP_1003J1_66_5789_n71 ) 
    , .SO ( DP_OP_1003J1_66_5789_n72 ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U44 (.A ( n1610 ) 
    , .B ( DP_OP_1003J1_66_5789_n69 ) , .CI ( DP_OP_1003J1_66_5789_n66 ) 
    , .CO ( DP_OP_1003J1_66_5789_n63 ) , .S ( DP_OP_1003J1_66_5789_n64 ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U45 (.A ( partial_3_L[12] ) 
    , .B ( partial_3_L[4] ) , .CI ( n1608 ) , .CO ( DP_OP_1003J1_66_5789_n65 ) 
    , .S ( DP_OP_1003J1_66_5789_n66 ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U42 (.A ( n1609 ) 
    , .B ( DP_OP_1003J1_66_5789_n65 ) , .CI ( DP_OP_1003J1_66_5789_n62 ) 
    , .CO ( DP_OP_1003J1_66_5789_n59 ) , .S ( DP_OP_1003J1_66_5789_n60 ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U43 (.A ( partial_3_L[13] ) 
    , .B ( partial_3_L[5] ) , .CI ( n1607 ) , .CO ( DP_OP_1003J1_66_5789_n61 ) 
    , .S ( DP_OP_1003J1_66_5789_n62 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U31 (.A ( DP_OP_1002J1_65_247_n41 ) , .B ( n1575 ) 
    , .CI ( DP_OP_1002J1_65_247_n44 ) , .CO ( DP_OP_1002J1_65_247_n38 ) 
    , .S ( DP_OP_1002J1_65_247_n39 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U34 (.A ( DP_OP_1002J1_65_247_n52 ) 
    , .B ( DP_OP_1002J1_65_247_n47 ) , .CI ( DP_OP_1002J1_65_247_n50 ) 
    , .CO ( DP_OP_1002J1_65_247_n44 ) , .S ( DP_OP_1002J1_65_247_n45 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U37 (.A ( DP_OP_1002J1_65_247_n58 ) 
    , .B ( DP_OP_1002J1_65_247_n53 ) , .CI ( DP_OP_1002J1_65_247_n56 ) 
    , .CO ( DP_OP_1002J1_65_247_n50 ) , .S ( DP_OP_1002J1_65_247_n51 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U40 (.A ( DP_OP_1002J1_65_247_n64 ) 
    , .B ( DP_OP_1002J1_65_247_n59 ) , .CI ( DP_OP_1002J1_65_247_n62 ) 
    , .CO ( DP_OP_1002J1_65_247_n56 ) , .S ( DP_OP_1002J1_65_247_n57 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U42 (.A ( sos2_reg_entrada[17] ) 
    , .B ( sos2_reg_entrada[15] ) , .CI ( sos2_reg_entrada[10] ) 
    , .CO ( DP_OP_1002J1_65_247_n60 ) , .S ( DP_OP_1002J1_65_247_n61 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U32 (.A ( DP_OP_1002J1_65_247_n48 ) 
    , .B ( DP_OP_1002J1_65_247_n43 ) , .CI ( DP_OP_1002J1_65_247_n46 ) 
    , .CO ( DP_OP_1002J1_65_247_n40 ) , .S ( DP_OP_1002J1_65_247_n41 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U28 (.A ( sos2_reg_entrada[17] ) 
    , .B ( sos2_reg_entrada[15] ) , .CI ( DP_OP_1002J1_65_247_n36 ) 
    , .CO ( DP_OP_1002J1_65_247_n32 ) , .S ( DP_OP_1002J1_65_247_n33 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U129 (.A ( DP_OP_1002J1_65_247_n184 ) 
    , .B ( DP_OP_1002J1_65_247_n183 ) , .CI ( DP_OP_1002J1_65_247_n164 ) 
    , .CO ( DP_OP_1002J1_65_247_n163 ) , .S ( DP_OP_1002J1_65_247_n273 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U9 (.A ( n1569 ) , .B ( DP_OP_1002J1_65_247_n23 ) 
    , .CI ( DP_OP_1002J1_65_247_n9 ) , .CO ( DP_OP_1002J1_65_247_n8 ) 
    , .S ( coeficiente_b12_H_v_out[11] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U11 (.A ( n1571 ) , .B ( DP_OP_1002J1_65_247_n27 ) 
    , .CI ( DP_OP_1002J1_65_247_n11 ) , .CO ( DP_OP_1002J1_65_247_n10 ) 
    , .S ( coeficiente_b12_H_v_out[9] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U14 (.A ( n1574 ) , .B ( DP_OP_1002J1_65_247_n39 ) 
    , .CI ( DP_OP_1002J1_65_247_n14 ) , .CO ( DP_OP_1002J1_65_247_n13 ) 
    , .S ( coeficiente_b12_H_v_out[6] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U16 (.A ( n1576 ) , .B ( DP_OP_1002J1_65_247_n51 ) 
    , .CI ( DP_OP_1002J1_65_247_n16 ) , .CO ( DP_OP_1002J1_65_247_n15 ) 
    , .S ( coeficiente_b12_H_v_out[4] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U17 (.A ( n1577 ) , .B ( DP_OP_1002J1_65_247_n57 ) 
    , .CI ( DP_OP_1002J1_65_247_n17 ) , .CO ( DP_OP_1002J1_65_247_n16 ) 
    , .S ( coeficiente_b12_H_v_out[3] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U25 (.A ( DP_OP_1002J1_65_247_n29 ) , .B ( n1572 ) 
    , .CI ( DP_OP_1002J1_65_247_n30 ) , .CO ( DP_OP_1002J1_65_247_n26 ) 
    , .S ( DP_OP_1002J1_65_247_n27 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U27 (.A ( DP_OP_1002J1_65_247_n33 ) , .B ( n1573 ) 
    , .CI ( DP_OP_1002J1_65_247_n34 ) , .CO ( DP_OP_1002J1_65_247_n30 ) 
    , .S ( DP_OP_1002J1_65_247_n31 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U29 (.A ( DP_OP_1002J1_65_247_n37 ) 
    , .B ( DP_OP_1002J1_65_247_n40 ) , .CI ( DP_OP_1002J1_65_247_n38 ) 
    , .CO ( DP_OP_1002J1_65_247_n34 ) , .S ( DP_OP_1002J1_65_247_n35 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U80 (.A ( n1580 ) , .B ( DP_OP_1002J1_65_247_n267 ) 
    , .CI ( DP_OP_1002J1_65_247_n106 ) , .CO ( DP_OP_1002J1_65_247_n105 ) 
    , .S ( coeficiente_b12_L_v_out[11] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U81 (.A ( DP_OP_1002J1_65_247_n130 ) 
    , .B ( DP_OP_1002J1_65_247_n266 ) , .CI ( DP_OP_1002J1_65_247_n107 ) 
    , .CO ( DP_OP_1002J1_65_247_n106 ) , .S ( coeficiente_b12_L_v_out[10] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U3 (.A ( n1564 ) , .B ( DP_OP_1002J1_65_247_n273 ) 
    , .CI ( DP_OP_1002J1_65_247_n3 ) , .CO ( DP_OP_1002J1_65_247_n2 ) 
    , .S ( coeficiente_b12_H_v_out[17] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U4 (.A ( n1565 ) , .B ( DP_OP_1002J1_65_247_n272 ) 
    , .CI ( DP_OP_1002J1_65_247_n4 ) , .CO ( DP_OP_1002J1_65_247_n3 ) 
    , .S ( coeficiente_b12_H_v_out[16] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U5 (.A ( n1566 ) , .B ( DP_OP_1002J1_65_247_n271 ) 
    , .CI ( DP_OP_1002J1_65_247_n5 ) , .CO ( DP_OP_1002J1_65_247_n4 ) 
    , .S ( coeficiente_b12_H_v_out[15] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U6 (.A ( n1567 ) , .B ( DP_OP_1002J1_65_247_n270 ) 
    , .CI ( DP_OP_1002J1_65_247_n6 ) , .CO ( DP_OP_1002J1_65_247_n5 ) 
    , .S ( coeficiente_b12_H_v_out[14] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U7 (.A ( n1568 ) , .B ( DP_OP_1002J1_65_247_n269 ) 
    , .CI ( DP_OP_1002J1_65_247_n7 ) , .CO ( DP_OP_1002J1_65_247_n6 ) 
    , .S ( coeficiente_b12_H_v_out[13] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U8 (.A ( DP_OP_1002J1_65_247_n22 ) 
    , .B ( DP_OP_1002J1_65_247_n268 ) , .CI ( DP_OP_1002J1_65_247_n8 ) 
    , .CO ( DP_OP_1002J1_65_247_n7 ) , .S ( coeficiente_b12_H_v_out[12] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U45 (.A ( sos2_reg_entrada[16] ) 
    , .B ( sos2_reg_entrada[14] ) , .CI ( sos2_reg_entrada[9] ) 
    , .CO ( DP_OP_1002J1_65_247_n66 ) , .S ( DP_OP_1002J1_65_247_n67 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U30 (.A ( sos2_reg_entrada[16] ) 
    , .B ( sos2_reg_entrada[14] ) , .CI ( DP_OP_1002J1_65_247_n42 ) 
    , .CO ( DP_OP_1002J1_65_247_n36 ) , .S ( DP_OP_1002J1_65_247_n37 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U133 (.A ( DP_OP_1002J1_65_247_n192 ) 
    , .B ( DP_OP_1002J1_65_247_n191 ) , .CI ( DP_OP_1002J1_65_247_n168 ) 
    , .CO ( DP_OP_1002J1_65_247_n167 ) , .S ( DP_OP_1002J1_65_247_n269 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U82 (.A ( DP_OP_1002J1_65_247_n132 ) 
    , .B ( DP_OP_1002J1_65_247_n265 ) , .CI ( DP_OP_1002J1_65_247_n108 ) 
    , .CO ( DP_OP_1002J1_65_247_n107 ) , .S ( coeficiente_b12_L_v_out[9] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U83 (.A ( DP_OP_1002J1_65_247_n134 ) 
    , .B ( DP_OP_1002J1_65_247_n264 ) , .CI ( DP_OP_1002J1_65_247_n109 ) 
    , .CO ( DP_OP_1002J1_65_247_n108 ) , .S ( coeficiente_b12_L_v_out[8] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U84 (.A ( DP_OP_1002J1_65_247_n136 ) 
    , .B ( DP_OP_1002J1_65_247_n263 ) , .CI ( DP_OP_1002J1_65_247_n110 ) 
    , .CO ( DP_OP_1002J1_65_247_n109 ) , .S ( coeficiente_b12_L_v_out[7] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U85 (.A ( DP_OP_1002J1_65_247_n138 ) 
    , .B ( DP_OP_1002J1_65_247_n262 ) , .CI ( DP_OP_1002J1_65_247_n111 ) 
    , .CO ( DP_OP_1002J1_65_247_n110 ) , .S ( coeficiente_b12_L_v_out[6] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U108 (.A ( sos2_reg_entrada[17] ) , .B ( n1585 ) 
    , .CI ( DP_OP_1002J1_65_247_n139 ) , .CO ( DP_OP_1002J1_65_247_n137 ) 
    , .S ( DP_OP_1002J1_65_247_n138 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U19 (.A ( DP_OP_1002J1_65_247_n19 ) , .B ( n1579 ) 
    , .CI ( DP_OP_1002J1_65_247_n69 ) , .CO ( DP_OP_1002J1_65_247_n18 ) 
    , .S ( coeficiente_b12_H_v_out[1] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U46 (.A ( DP_OP_1002J1_65_247_n73 ) , .B ( n1589 ) 
    , .CI ( DP_OP_1002J1_65_247_n71 ) , .CO ( DP_OP_1002J1_65_247_n68 ) 
    , .S ( DP_OP_1002J1_65_247_n69 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U47 (.A ( sos2_reg_entrada[15] ) 
    , .B ( sos2_reg_entrada[10] ) , .CI ( DP_OP_1002J1_65_247_n74 ) 
    , .CO ( DP_OP_1002J1_65_247_n70 ) , .S ( DP_OP_1002J1_65_247_n71 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U134 (.A ( DP_OP_1002J1_65_247_n194 ) 
    , .B ( DP_OP_1002J1_65_247_n193 ) , .CI ( DP_OP_1002J1_65_247_n169 ) 
    , .CO ( DP_OP_1002J1_65_247_n168 ) , .S ( DP_OP_1002J1_65_247_n268 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U86 (.A ( DP_OP_1002J1_65_247_n140 ) 
    , .B ( DP_OP_1002J1_65_247_n261 ) , .CI ( DP_OP_1002J1_65_247_n112 ) 
    , .CO ( DP_OP_1002J1_65_247_n111 ) , .S ( coeficiente_b12_L_v_out[5] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U109 (.A ( sos2_reg_entrada[16] ) , .B ( n1584 ) 
    , .CI ( DP_OP_1002J1_65_247_n141 ) , .CO ( DP_OP_1002J1_65_247_n139 ) 
    , .S ( DP_OP_1002J1_65_247_n140 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U18 (.A ( n1578 ) , .B ( DP_OP_1002J1_65_247_n63 ) 
    , .CI ( DP_OP_1002J1_65_247_n18 ) , .CO ( DP_OP_1002J1_65_247_n17 ) 
    , .S ( coeficiente_b12_H_v_out[2] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U43 (.A ( DP_OP_1002J1_65_247_n70 ) 
    , .B ( DP_OP_1002J1_65_247_n65 ) , .CI ( DP_OP_1002J1_65_247_n68 ) 
    , .CO ( DP_OP_1002J1_65_247_n62 ) , .S ( DP_OP_1002J1_65_247_n63 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U112 (.A ( sos2_reg_entrada[13] ) , .B ( n1581 ) 
    , .CI ( DP_OP_1002J1_65_247_n147 ) , .CO ( DP_OP_1002J1_65_247_n145 ) 
    , .S ( DP_OP_1002J1_65_247_n146 ) ) ;
HADDX1 DP_OP_1002J1_65_247_U48 (.B0 ( sos2_reg_entrada[8] ) 
    , .A0 ( sos2_reg_entrada[13] ) , .C1 ( DP_OP_1002J1_65_247_n72 ) 
    , .SO ( DP_OP_1002J1_65_247_n73 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U136 (.A ( DP_OP_1002J1_65_247_n198 ) 
    , .B ( DP_OP_1002J1_65_247_n197 ) , .CI ( DP_OP_1002J1_65_247_n171 ) 
    , .CO ( DP_OP_1002J1_65_247_n170 ) , .S ( DP_OP_1002J1_65_247_n266 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U88 (.A ( DP_OP_1002J1_65_247_n144 ) 
    , .B ( DP_OP_1002J1_65_247_n259 ) , .CI ( DP_OP_1002J1_65_247_n114 ) 
    , .CO ( DP_OP_1002J1_65_247_n113 ) , .S ( coeficiente_b12_L_v_out[3] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U111 (.A ( sos2_reg_entrada[14] ) , .B ( n1582 ) 
    , .CI ( DP_OP_1002J1_65_247_n145 ) , .CO ( DP_OP_1002J1_65_247_n143 ) 
    , .S ( DP_OP_1002J1_65_247_n144 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U20 (.A ( sos2_reg_entrada[14] ) 
    , .B ( DP_OP_1002J1_65_247_n75 ) , .CI ( DP_OP_1002J1_65_247_n256 ) 
    , .CO ( DP_OP_1002J1_65_247_n19 ) , .S ( coeficiente_b12_H_v_out[0] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U135 (.A ( DP_OP_1002J1_65_247_n196 ) 
    , .B ( DP_OP_1002J1_65_247_n195 ) , .CI ( DP_OP_1002J1_65_247_n170 ) 
    , .CO ( DP_OP_1002J1_65_247_n169 ) , .S ( DP_OP_1002J1_65_247_n267 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U87 (.A ( DP_OP_1002J1_65_247_n142 ) 
    , .B ( DP_OP_1002J1_65_247_n260 ) , .CI ( DP_OP_1002J1_65_247_n113 ) 
    , .CO ( DP_OP_1002J1_65_247_n112 ) , .S ( coeficiente_b12_L_v_out[4] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U140 (.A ( DP_OP_1002J1_65_247_n206 ) 
    , .B ( DP_OP_1002J1_65_247_n205 ) , .CI ( DP_OP_1002J1_65_247_n175 ) 
    , .CO ( DP_OP_1002J1_65_247_n174 ) , .S ( DP_OP_1002J1_65_247_n262 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U139 (.A ( DP_OP_1002J1_65_247_n204 ) 
    , .B ( DP_OP_1002J1_65_247_n203 ) , .CI ( DP_OP_1002J1_65_247_n174 ) 
    , .CO ( DP_OP_1002J1_65_247_n173 ) , .S ( DP_OP_1002J1_65_247_n263 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U91 (.A ( sos2_reg_entrada[11] ) 
    , .B ( sos2_reg_entrada[8] ) , .CI ( DP_OP_1002J1_65_247_n256 ) 
    , .CO ( DP_OP_1002J1_65_247_n116 ) , .S ( coeficiente_b12_L_v_out[0] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U138 (.A ( DP_OP_1002J1_65_247_n202 ) 
    , .B ( DP_OP_1002J1_65_247_n201 ) , .CI ( DP_OP_1002J1_65_247_n173 ) 
    , .CO ( DP_OP_1002J1_65_247_n172 ) , .S ( DP_OP_1002J1_65_247_n264 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U90 (.A ( DP_OP_1002J1_65_247_n148 ) 
    , .B ( DP_OP_1002J1_65_247_n116 ) , .CI ( DP_OP_1002J1_65_247_n257 ) 
    , .CO ( DP_OP_1002J1_65_247_n115 ) , .S ( coeficiente_b12_L_v_out[1] ) ) ;
FADDX1 DP_OP_1002J1_65_247_U113 (.A ( sos2_reg_entrada[12] ) , .B ( n1597 ) 
    , .CI ( n1596 ) , .CO ( DP_OP_1002J1_65_247_n147 ) 
    , .S ( DP_OP_1002J1_65_247_n148 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U137 (.A ( DP_OP_1002J1_65_247_n200 ) 
    , .B ( DP_OP_1002J1_65_247_n199 ) , .CI ( DP_OP_1002J1_65_247_n172 ) 
    , .CO ( DP_OP_1002J1_65_247_n171 ) , .S ( DP_OP_1002J1_65_247_n265 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U89 (.A ( DP_OP_1002J1_65_247_n146 ) 
    , .B ( DP_OP_1002J1_65_247_n258 ) , .CI ( DP_OP_1002J1_65_247_n115 ) 
    , .CO ( DP_OP_1002J1_65_247_n114 ) , .S ( coeficiente_b12_L_v_out[2] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U258 (.A ( in_reg_salida_v[17] ) , .B ( n1539 ) 
    , .CI ( coeficiente_a22_in[18] ) , .CO ( DP_OP_1001J1_64_4995_n336 ) 
    , .S ( DP_OP_1001J1_64_4995_n337 ) ) ;
HADDX1 DP_OP_1002J1_65_247_U146 (.B0 ( n1591 ) , .A0 ( n1590 ) 
    , .C1 ( DP_OP_1002J1_65_247_n180 ) , .SO ( DP_OP_1002J1_65_247_n256 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U145 (.A ( n1592 ) 
    , .B ( DP_OP_1002J1_65_247_n180 ) , .CI ( DP_OP_1002J1_65_247_n215 ) 
    , .CO ( DP_OP_1002J1_65_247_n179 ) , .S ( DP_OP_1002J1_65_247_n257 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U144 (.A ( DP_OP_1002J1_65_247_n214 ) 
    , .B ( DP_OP_1002J1_65_247_n213 ) , .CI ( DP_OP_1002J1_65_247_n179 ) 
    , .CO ( DP_OP_1002J1_65_247_n178 ) , .S ( DP_OP_1002J1_65_247_n258 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U143 (.A ( DP_OP_1002J1_65_247_n212 ) 
    , .B ( DP_OP_1002J1_65_247_n211 ) , .CI ( DP_OP_1002J1_65_247_n178 ) 
    , .CO ( DP_OP_1002J1_65_247_n177 ) , .S ( DP_OP_1002J1_65_247_n259 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U162 (.A ( sos2_reg_entrada[2] ) , .B ( n1592 ) 
    , .CI ( n1594 ) , .CO ( DP_OP_1002J1_65_247_n210 ) 
    , .S ( DP_OP_1002J1_65_247_n211 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U142 (.A ( DP_OP_1002J1_65_247_n210 ) 
    , .B ( DP_OP_1002J1_65_247_n209 ) , .CI ( DP_OP_1002J1_65_247_n177 ) 
    , .CO ( DP_OP_1002J1_65_247_n176 ) , .S ( DP_OP_1002J1_65_247_n260 ) ) ;
FADDX1 DP_OP_1002J1_65_247_U141 (.A ( DP_OP_1002J1_65_247_n208 ) 
    , .B ( DP_OP_1002J1_65_247_n207 ) , .CI ( DP_OP_1002J1_65_247_n176 ) 
    , .CO ( DP_OP_1002J1_65_247_n175 ) , .S ( DP_OP_1002J1_65_247_n261 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U285 (.A ( DP_OP_1001J1_64_4995_n406 ) 
    , .B ( DP_OP_1001J1_64_4995_n395 ) , .CI ( DP_OP_1001J1_64_4995_n404 ) 
    , .CO ( DP_OP_1001J1_64_4995_n390 ) , .S ( DP_OP_1001J1_64_4995_n391 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U292 (.A ( DP_OP_1001J1_64_4995_n420 ) 
    , .B ( DP_OP_1001J1_64_4995_n411 ) , .CI ( DP_OP_1001J1_64_4995_n409 ) 
    , .CO ( DP_OP_1001J1_64_4995_n404 ) , .S ( DP_OP_1001J1_64_4995_n405 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U275 (.A ( DP_OP_1001J1_64_4995_n375 ) 
    , .B ( DP_OP_1001J1_64_4995_n380 ) , .CI ( DP_OP_1001J1_64_4995_n373 ) 
    , .CO ( DP_OP_1001J1_64_4995_n370 ) , .S ( DP_OP_1001J1_64_4995_n371 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U280 (.A ( DP_OP_1001J1_64_4995_n385 ) 
    , .B ( DP_OP_1001J1_64_4995_n394 ) , .CI ( DP_OP_1001J1_64_4995_n392 ) 
    , .CO ( DP_OP_1001J1_64_4995_n380 ) , .S ( DP_OP_1001J1_64_4995_n381 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U287 (.A ( coeficiente_a22_in[18] ) 
    , .B ( sos2_reg_entrada[18] ) , .CI ( DP_OP_1001J1_64_4995_n410 ) 
    , .CO ( DP_OP_1001J1_64_4995_n394 ) , .S ( DP_OP_1001J1_64_4995_n395 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U265 (.A ( DP_OP_1001J1_64_4995_n355 ) 
    , .B ( DP_OP_1001J1_64_4995_n358 ) , .CI ( DP_OP_1001J1_64_4995_n353 ) 
    , .CO ( DP_OP_1001J1_64_4995_n350 ) , .S ( DP_OP_1001J1_64_4995_n351 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U263 (.A ( DP_OP_1001J1_64_4995_n354 ) 
    , .B ( DP_OP_1001J1_64_4995_n349 ) , .CI ( DP_OP_1001J1_64_4995_n352 ) 
    , .CO ( DP_OP_1001J1_64_4995_n346 ) , .S ( DP_OP_1001J1_64_4995_n347 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U266 (.A ( n1534 ) , .B ( n1540 ) 
    , .CI ( DP_OP_1001J1_64_4995_n360 ) , .CO ( DP_OP_1001J1_64_4995_n352 ) 
    , .S ( DP_OP_1001J1_64_4995_n353 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U249 (.A ( DP_OP_1001J1_64_4995_n412 ) 
    , .B ( DP_OP_1001J1_64_4995_n401 ) , .CI ( DP_OP_1001J1_64_4995_n328 ) 
    , .CO ( DP_OP_1001J1_64_4995_n327 ) , .S ( partial_1[6] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U250 (.A ( DP_OP_1001J1_64_4995_n426 ) 
    , .B ( DP_OP_1001J1_64_4995_n413 ) , .CI ( DP_OP_1001J1_64_4995_n329 ) 
    , .CO ( DP_OP_1001J1_64_4995_n328 ) , .S ( partial_1[5] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U296 (.A ( DP_OP_1001J1_64_4995_n417 ) 
    , .B ( DP_OP_1001J1_64_4995_n428 ) , .CI ( DP_OP_1001J1_64_4995_n415 ) 
    , .CO ( DP_OP_1001J1_64_4995_n412 ) , .S ( DP_OP_1001J1_64_4995_n413 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U290 (.A ( DP_OP_1001J1_64_4995_n405 ) 
    , .B ( DP_OP_1001J1_64_4995_n414 ) , .CI ( DP_OP_1001J1_64_4995_n403 ) 
    , .CO ( DP_OP_1001J1_64_4995_n400 ) , .S ( DP_OP_1001J1_64_4995_n401 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U284 (.A ( DP_OP_1001J1_64_4995_n393 ) 
    , .B ( DP_OP_1001J1_64_4995_n402 ) , .CI ( DP_OP_1001J1_64_4995_n391 ) 
    , .CO ( DP_OP_1001J1_64_4995_n388 ) , .S ( DP_OP_1001J1_64_4995_n389 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U291 (.A ( DP_OP_1001J1_64_4995_n418 ) 
    , .B ( DP_OP_1001J1_64_4995_n407 ) , .CI ( DP_OP_1001J1_64_4995_n416 ) 
    , .CO ( DP_OP_1001J1_64_4995_n402 ) , .S ( DP_OP_1001J1_64_4995_n403 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U298 (.A ( DP_OP_1001J1_64_4995_n425 ) 
    , .B ( DP_OP_1001J1_64_4995_n423 ) , .CI ( DP_OP_1001J1_64_4995_n421 ) 
    , .CO ( DP_OP_1001J1_64_4995_n416 ) , .S ( DP_OP_1001J1_64_4995_n417 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U279 (.A ( DP_OP_1001J1_64_4995_n383 ) 
    , .B ( DP_OP_1001J1_64_4995_n390 ) , .CI ( DP_OP_1001J1_64_4995_n381 ) 
    , .CO ( DP_OP_1001J1_64_4995_n378 ) , .S ( DP_OP_1001J1_64_4995_n379 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U34 (.A ( DP_OP_1001J1_64_4995_n83 ) 
    , .B ( DP_OP_1001J1_64_4995_n558 ) , .CI ( DP_OP_1001J1_64_4995_n33 ) 
    , .CO ( DP_OP_1001J1_64_4995_n32 ) , .S ( partial_2_H[8] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U35 (.A ( DP_OP_1001J1_64_4995_n87 ) 
    , .B ( DP_OP_1001J1_64_4995_n557 ) , .CI ( DP_OP_1001J1_64_4995_n34 ) 
    , .CO ( DP_OP_1001J1_64_4995_n33 ) , .S ( partial_2_H[7] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U36 (.A ( DP_OP_1001J1_64_4995_n93 ) 
    , .B ( DP_OP_1001J1_64_4995_n556 ) , .CI ( DP_OP_1001J1_64_4995_n35 ) 
    , .CO ( DP_OP_1001J1_64_4995_n34 ) , .S ( partial_2_H[6] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U37 (.A ( DP_OP_1001J1_64_4995_n99 ) 
    , .B ( DP_OP_1001J1_64_4995_n555 ) , .CI ( DP_OP_1001J1_64_4995_n36 ) 
    , .CO ( DP_OP_1001J1_64_4995_n35 ) , .S ( partial_2_H[5] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U228 (.A ( coeficiente_a22_in[7] ) 
    , .B ( partial_1[7] ) , .CI ( DP_OP_1001J1_64_4995_n308 ) 
    , .CO ( DP_OP_1001J1_64_4995_n307 ) , .S ( DP_OP_1001J1_64_4995_n557 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U229 (.A ( coeficiente_a22_in[6] ) 
    , .B ( partial_1[6] ) , .CI ( DP_OP_1001J1_64_4995_n309 ) 
    , .CO ( DP_OP_1001J1_64_4995_n308 ) , .S ( DP_OP_1001J1_64_4995_n556 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U230 (.A ( coeficiente_a22_in[5] ) 
    , .B ( partial_1[5] ) , .CI ( DP_OP_1001J1_64_4995_n310 ) 
    , .CO ( DP_OP_1001J1_64_4995_n309 ) , .S ( DP_OP_1001J1_64_4995_n555 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U248 (.A ( DP_OP_1001J1_64_4995_n400 ) 
    , .B ( DP_OP_1001J1_64_4995_n389 ) , .CI ( DP_OP_1001J1_64_4995_n327 ) 
    , .CO ( DP_OP_1001J1_64_4995_n326 ) , .S ( partial_1[7] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U10 (.A ( coeficiente_b11_H_v_out[11] ) 
    , .B ( partial_2_H[11] ) , .CI ( DP_OP_1001J1_64_4995_n10 ) 
    , .CO ( DP_OP_1001J1_64_4995_n9 ) , .S ( partial_3_H[11] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U11 (.A ( coeficiente_b11_H_v_out[10] ) 
    , .B ( partial_2_H[10] ) , .CI ( DP_OP_1001J1_64_4995_n11 ) 
    , .CO ( DP_OP_1001J1_64_4995_n10 ) , .S ( partial_3_H[10] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U12 (.A ( coeficiente_b11_H_v_out[9] ) 
    , .B ( partial_2_H[9] ) , .CI ( DP_OP_1001J1_64_4995_n12 ) 
    , .CO ( DP_OP_1001J1_64_4995_n11 ) , .S ( partial_3_H[9] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U13 (.A ( coeficiente_b11_H_v_out[8] ) 
    , .B ( partial_2_H[8] ) , .CI ( DP_OP_1001J1_64_4995_n13 ) 
    , .CO ( DP_OP_1001J1_64_4995_n12 ) , .S ( partial_3_H[8] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U14 (.A ( coeficiente_b11_H_v_out[7] ) 
    , .B ( partial_2_H[7] ) , .CI ( DP_OP_1001J1_64_4995_n14 ) 
    , .CO ( DP_OP_1001J1_64_4995_n13 ) , .S ( partial_3_H[7] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U15 (.A ( coeficiente_b11_H_v_out[6] ) 
    , .B ( partial_2_H[6] ) , .CI ( DP_OP_1001J1_64_4995_n15 ) 
    , .CO ( DP_OP_1001J1_64_4995_n14 ) , .S ( partial_3_H[6] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U16 (.A ( coeficiente_b11_H_v_out[5] ) 
    , .B ( partial_2_H[5] ) , .CI ( DP_OP_1001J1_64_4995_n16 ) 
    , .CO ( DP_OP_1001J1_64_4995_n15 ) , .S ( partial_3_H[5] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U32 (.A ( DP_OP_1001J1_64_4995_n75 ) 
    , .B ( DP_OP_1001J1_64_4995_n560 ) , .CI ( DP_OP_1001J1_64_4995_n31 ) 
    , .CO ( DP_OP_1001J1_64_4995_n30 ) , .S ( partial_2_H[10] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U121 (.A ( coeficiente_b11_L_v_out[7] ) 
    , .B ( partial_2_L[7] ) , .CI ( DP_OP_1001J1_64_4995_n161 ) 
    , .CO ( DP_OP_1001J1_64_4995_n160 ) , .S ( partial_3_L[7] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U122 (.A ( coeficiente_b11_L_v_out[6] ) 
    , .B ( partial_2_L[6] ) , .CI ( DP_OP_1001J1_64_4995_n162 ) 
    , .CO ( DP_OP_1001J1_64_4995_n161 ) , .S ( partial_3_L[6] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U123 (.A ( coeficiente_b11_L_v_out[5] ) 
    , .B ( partial_2_L[5] ) , .CI ( DP_OP_1001J1_64_4995_n163 ) 
    , .CO ( DP_OP_1001J1_64_4995_n162 ) , .S ( partial_3_L[5] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U142 (.A ( DP_OP_1001J1_64_4995_n234 ) 
    , .B ( DP_OP_1001J1_64_4995_n557 ) , .CI ( DP_OP_1001J1_64_4995_n181 ) 
    , .CO ( DP_OP_1001J1_64_4995_n180 ) , .S ( partial_2_L[7] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U143 (.A ( DP_OP_1001J1_64_4995_n240 ) 
    , .B ( DP_OP_1001J1_64_4995_n556 ) , .CI ( DP_OP_1001J1_64_4995_n182 ) 
    , .CO ( DP_OP_1001J1_64_4995_n181 ) , .S ( partial_2_L[6] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U144 (.A ( DP_OP_1001J1_64_4995_n246 ) 
    , .B ( DP_OP_1001J1_64_4995_n555 ) , .CI ( DP_OP_1001J1_64_4995_n183 ) 
    , .CO ( DP_OP_1001J1_64_4995_n182 ) , .S ( partial_2_L[5] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U6 (.A ( coeficiente_b11_H_v_out[15] ) 
    , .B ( partial_2_H[15] ) , .CI ( DP_OP_1001J1_64_4995_n6 ) 
    , .CO ( DP_OP_1001J1_64_4995_n5 ) , .S ( partial_3_H[15] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U9 (.A ( coeficiente_b11_H_v_out[12] ) 
    , .B ( partial_2_H[12] ) , .CI ( DP_OP_1001J1_64_4995_n9 ) 
    , .CO ( DP_OP_1001J1_64_4995_n8 ) , .S ( partial_3_H[12] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U111 (.A ( coeficiente_b11_L_v_out[17] ) 
    , .B ( partial_2_L[17] ) , .CI ( DP_OP_1001J1_64_4995_n151 ) 
    , .CO ( DP_OP_1001J1_64_4995_n150 ) , .S ( partial_3_L[17] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U112 (.A ( coeficiente_b11_L_v_out[16] ) 
    , .B ( partial_2_L[16] ) , .CI ( DP_OP_1001J1_64_4995_n152 ) 
    , .CO ( DP_OP_1001J1_64_4995_n151 ) , .S ( partial_3_L[16] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U113 (.A ( coeficiente_b11_L_v_out[15] ) 
    , .B ( partial_2_L[15] ) , .CI ( DP_OP_1001J1_64_4995_n153 ) 
    , .CO ( DP_OP_1001J1_64_4995_n152 ) , .S ( partial_3_L[15] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U114 (.A ( coeficiente_b11_L_v_out[14] ) 
    , .B ( partial_2_L[14] ) , .CI ( DP_OP_1001J1_64_4995_n154 ) 
    , .CO ( DP_OP_1001J1_64_4995_n153 ) , .S ( partial_3_L[14] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U115 (.A ( coeficiente_b11_L_v_out[13] ) 
    , .B ( partial_2_L[13] ) , .CI ( DP_OP_1001J1_64_4995_n155 ) 
    , .CO ( DP_OP_1001J1_64_4995_n154 ) , .S ( partial_3_L[13] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U116 (.A ( coeficiente_b11_L_v_out[12] ) 
    , .B ( partial_2_L[12] ) , .CI ( DP_OP_1001J1_64_4995_n156 ) 
    , .CO ( DP_OP_1001J1_64_4995_n155 ) , .S ( partial_3_L[12] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U119 (.A ( coeficiente_b11_L_v_out[9] ) 
    , .B ( partial_2_L[9] ) , .CI ( DP_OP_1001J1_64_4995_n159 ) 
    , .CO ( DP_OP_1001J1_64_4995_n158 ) , .S ( partial_3_L[9] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U120 (.A ( coeficiente_b11_L_v_out[8] ) 
    , .B ( partial_2_L[8] ) , .CI ( DP_OP_1001J1_64_4995_n160 ) 
    , .CO ( DP_OP_1001J1_64_4995_n159 ) , .S ( partial_3_L[8] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U251 (.A ( DP_OP_1001J1_64_4995_n440 ) 
    , .B ( DP_OP_1001J1_64_4995_n427 ) , .CI ( DP_OP_1001J1_64_4995_n330 ) 
    , .CO ( DP_OP_1001J1_64_4995_n329 ) , .S ( partial_1[4] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U303 (.A ( DP_OP_1001J1_64_4995_n431 ) 
    , .B ( DP_OP_1001J1_64_4995_n442 ) , .CI ( DP_OP_1001J1_64_4995_n429 ) 
    , .CO ( DP_OP_1001J1_64_4995_n426 ) , .S ( DP_OP_1001J1_64_4995_n427 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U297 (.A ( DP_OP_1001J1_64_4995_n432 ) 
    , .B ( DP_OP_1001J1_64_4995_n430 ) , .CI ( DP_OP_1001J1_64_4995_n419 ) 
    , .CO ( DP_OP_1001J1_64_4995_n414 ) , .S ( DP_OP_1001J1_64_4995_n415 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U305 (.A ( DP_OP_1001J1_64_4995_n439 ) 
    , .B ( DP_OP_1001J1_64_4995_n437 ) , .CI ( DP_OP_1001J1_64_4995_n435 ) 
    , .CO ( DP_OP_1001J1_64_4995_n430 ) , .S ( DP_OP_1001J1_64_4995_n431 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U299 (.A ( DP_OP_1001J1_64_4995_n438 ) 
    , .B ( DP_OP_1001J1_64_4995_n436 ) , .CI ( DP_OP_1001J1_64_4995_n434 ) 
    , .CO ( DP_OP_1001J1_64_4995_n418 ) , .S ( DP_OP_1001J1_64_4995_n419 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U309 (.A ( in_reg_salida_v[4] ) 
    , .B ( coeficiente_a22_in[8] ) , .CI ( coeficiente_a22_in[17] ) 
    , .CO ( DP_OP_1001J1_64_4995_n438 ) , .S ( DP_OP_1001J1_64_4995_n439 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U268 (.A ( DP_OP_1001J1_64_4995_n361 ) 
    , .B ( DP_OP_1001J1_64_4995_n364 ) , .CI ( DP_OP_1001J1_64_4995_n359 ) 
    , .CO ( DP_OP_1001J1_64_4995_n356 ) , .S ( DP_OP_1001J1_64_4995_n357 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U286 (.A ( DP_OP_1001J1_64_4995_n408 ) 
    , .B ( DP_OP_1001J1_64_4995_n399 ) , .CI ( DP_OP_1001J1_64_4995_n397 ) 
    , .CO ( DP_OP_1001J1_64_4995_n392 ) , .S ( DP_OP_1001J1_64_4995_n393 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U272 (.A ( DP_OP_1001J1_64_4995_n376 ) 
    , .B ( DP_OP_1001J1_64_4995_n369 ) , .CI ( DP_OP_1001J1_64_4995_n367 ) 
    , .CO ( DP_OP_1001J1_64_4995_n364 ) , .S ( DP_OP_1001J1_64_4995_n365 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U274 (.A ( in_reg_salida_v[10] ) 
    , .B ( coeficiente_a22_in[14] ) , .CI ( coeficiente_a22_in[16] ) 
    , .CO ( DP_OP_1001J1_64_4995_n368 ) , .S ( DP_OP_1001J1_64_4995_n369 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U267 (.A ( in_reg_salida_v[12] ) 
    , .B ( coeficiente_a22_in[16] ) , .CI ( n1535 ) 
    , .CO ( DP_OP_1001J1_64_4995_n354 ) , .S ( DP_OP_1001J1_64_4995_n355 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U124 (.A ( coeficiente_b11_L_v_out[4] ) 
    , .B ( DP_OP_1001J1_64_4995_n164 ) , .CI ( partial_2_L[4] ) 
    , .CO ( DP_OP_1001J1_64_4995_n163 ) , .S ( partial_3_L[4] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U145 (.A ( DP_OP_1001J1_64_4995_n252 ) 
    , .B ( DP_OP_1001J1_64_4995_n554 ) , .CI ( DP_OP_1001J1_64_4995_n184 ) 
    , .CO ( DP_OP_1001J1_64_4995_n183 ) , .S ( partial_2_L[4] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U17 (.A ( coeficiente_b11_H_v_out[4] ) 
    , .B ( DP_OP_1001J1_64_4995_n17 ) , .CI ( partial_2_H[4] ) 
    , .CO ( DP_OP_1001J1_64_4995_n16 ) , .S ( partial_3_H[4] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U38 (.A ( DP_OP_1001J1_64_4995_n105 ) 
    , .B ( DP_OP_1001J1_64_4995_n554 ) , .CI ( DP_OP_1001J1_64_4995_n37 ) 
    , .CO ( DP_OP_1001J1_64_4995_n36 ) , .S ( partial_2_H[4] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U231 (.A ( coeficiente_a22_in[4] ) 
    , .B ( partial_1[4] ) , .CI ( DP_OP_1001J1_64_4995_n311 ) 
    , .CO ( DP_OP_1001J1_64_4995_n310 ) , .S ( DP_OP_1001J1_64_4995_n554 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U125 (.A ( coeficiente_b11_L_v_out[3] ) 
    , .B ( DP_OP_1001J1_64_4995_n165 ) , .CI ( partial_2_L[3] ) 
    , .CO ( DP_OP_1001J1_64_4995_n164 ) , .S ( partial_3_L[3] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U18 (.A ( coeficiente_b11_H_v_out[3] ) 
    , .B ( DP_OP_1001J1_64_4995_n18 ) , .CI ( partial_2_H[3] ) 
    , .CO ( DP_OP_1001J1_64_4995_n17 ) , .S ( partial_3_H[3] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U310 (.A ( DP_OP_1001J1_64_4995_n445 ) 
    , .B ( DP_OP_1001J1_64_4995_n456 ) , .CI ( DP_OP_1001J1_64_4995_n443 ) 
    , .CO ( DP_OP_1001J1_64_4995_n440 ) , .S ( DP_OP_1001J1_64_4995_n441 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U304 (.A ( DP_OP_1001J1_64_4995_n446 ) 
    , .B ( DP_OP_1001J1_64_4995_n444 ) , .CI ( DP_OP_1001J1_64_4995_n433 ) 
    , .CO ( DP_OP_1001J1_64_4995_n428 ) , .S ( DP_OP_1001J1_64_4995_n429 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U312 (.A ( DP_OP_1001J1_64_4995_n453 ) 
    , .B ( DP_OP_1001J1_64_4995_n451 ) , .CI ( DP_OP_1001J1_64_4995_n449 ) 
    , .CO ( DP_OP_1001J1_64_4995_n444 ) , .S ( DP_OP_1001J1_64_4995_n445 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U306 (.A ( DP_OP_1001J1_64_4995_n452 ) 
    , .B ( DP_OP_1001J1_64_4995_n450 ) , .CI ( DP_OP_1001J1_64_4995_n448 ) 
    , .CO ( DP_OP_1001J1_64_4995_n432 ) , .S ( DP_OP_1001J1_64_4995_n433 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U316 (.A ( in_reg_salida_v[3] ) 
    , .B ( coeficiente_a22_in[7] ) , .CI ( coeficiente_a22_in[16] ) 
    , .CO ( DP_OP_1001J1_64_4995_n452 ) , .S ( DP_OP_1001J1_64_4995_n453 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U271 (.A ( DP_OP_1001J1_64_4995_n374 ) 
    , .B ( DP_OP_1001J1_64_4995_n372 ) , .CI ( DP_OP_1001J1_64_4995_n365 ) 
    , .CO ( DP_OP_1001J1_64_4995_n362 ) , .S ( DP_OP_1001J1_64_4995_n363 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U126 (.A ( coeficiente_b11_L_v_out[2] ) 
    , .B ( DP_OP_1001J1_64_4995_n166 ) , .CI ( partial_2_L[2] ) 
    , .CO ( DP_OP_1001J1_64_4995_n165 ) , .S ( partial_3_L[2] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U19 (.A ( coeficiente_b11_H_v_out[2] ) 
    , .B ( DP_OP_1001J1_64_4995_n19 ) , .CI ( partial_2_H[2] ) 
    , .CO ( DP_OP_1001J1_64_4995_n18 ) , .S ( partial_3_H[2] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U317 (.A ( DP_OP_1001J1_64_4995_n461 ) 
    , .B ( DP_OP_1001J1_64_4995_n459 ) , .CI ( DP_OP_1001J1_64_4995_n468 ) 
    , .CO ( DP_OP_1001J1_64_4995_n454 ) , .S ( DP_OP_1001J1_64_4995_n455 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U311 (.A ( DP_OP_1001J1_64_4995_n460 ) 
    , .B ( DP_OP_1001J1_64_4995_n458 ) , .CI ( DP_OP_1001J1_64_4995_n447 ) 
    , .CO ( DP_OP_1001J1_64_4995_n442 ) , .S ( DP_OP_1001J1_64_4995_n443 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U319 (.A ( DP_OP_1001J1_64_4995_n474 ) 
    , .B ( DP_OP_1001J1_64_4995_n467 ) , .CI ( DP_OP_1001J1_64_4995_n465 ) 
    , .CO ( DP_OP_1001J1_64_4995_n458 ) , .S ( DP_OP_1001J1_64_4995_n459 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U313 (.A ( DP_OP_1001J1_64_4995_n466 ) 
    , .B ( DP_OP_1001J1_64_4995_n464 ) , .CI ( DP_OP_1001J1_64_4995_n462 ) 
    , .CO ( DP_OP_1001J1_64_4995_n446 ) , .S ( DP_OP_1001J1_64_4995_n447 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U307 (.A ( n1537 ) , .B ( n1586 ) , .CI ( n1545 ) 
    , .CO ( DP_OP_1001J1_64_4995_n434 ) , .S ( DP_OP_1001J1_64_4995_n435 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U262 (.A ( in_reg_salida_v[14] ) , .B ( n1536 ) 
    , .CI ( n1537 ) , .CO ( DP_OP_1001J1_64_4995_n344 ) 
    , .S ( DP_OP_1001J1_64_4995_n345 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U327 (.A ( n1597 ) , .B ( n1534 ) 
    , .CI ( DP_OP_1001J1_64_4995_n484 ) , .CO ( DP_OP_1001J1_64_4995_n472 ) 
    , .S ( DP_OP_1001J1_64_4995_n473 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U289 (.A ( sos2_reg_entrada[15] ) 
    , .B ( coeficiente_a22_in[13] ) , .CI ( coeficiente_a22_in[11] ) 
    , .CO ( DP_OP_1001J1_64_4995_n398 ) , .S ( DP_OP_1001J1_64_4995_n399 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U325 (.A ( DP_OP_1001J1_64_4995_n477 ) 
    , .B ( DP_OP_1001J1_64_4995_n475 ) , .CI ( DP_OP_1001J1_64_4995_n473 ) 
    , .CO ( DP_OP_1001J1_64_4995_n468 ) , .S ( DP_OP_1001J1_64_4995_n469 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U281 (.A ( DP_OP_1001J1_64_4995_n398 ) 
    , .B ( DP_OP_1001J1_64_4995_n396 ) , .CI ( DP_OP_1001J1_64_4995_n387 ) 
    , .CO ( DP_OP_1001J1_64_4995_n382 ) , .S ( DP_OP_1001J1_64_4995_n383 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U283 (.A ( in_reg_salida_v[8] ) 
    , .B ( coeficiente_a22_in[14] ) , .CI ( coeficiente_a22_in[12] ) 
    , .CO ( DP_OP_1001J1_64_4995_n386 ) , .S ( DP_OP_1001J1_64_4995_n387 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U314 (.A ( n1536 ) , .B ( n1585 ) , .CI ( n1544 ) 
    , .CO ( DP_OP_1001J1_64_4995_n448 ) , .S ( DP_OP_1001J1_64_4995_n449 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U276 (.A ( DP_OP_1001J1_64_4995_n384 ) 
    , .B ( DP_OP_1001J1_64_4995_n377 ) , .CI ( DP_OP_1001J1_64_4995_n382 ) 
    , .CO ( DP_OP_1001J1_64_4995_n372 ) , .S ( DP_OP_1001J1_64_4995_n373 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U278 (.A ( sos2_reg_entrada[17] ) 
    , .B ( in_reg_salida_v[9] ) , .CI ( coeficiente_a22_in[15] ) 
    , .CO ( DP_OP_1001J1_64_4995_n376 ) , .S ( DP_OP_1001J1_64_4995_n377 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U293 (.A ( n1547 ) 
    , .B ( DP_OP_1001J1_64_4995_n424 ) , .CI ( DP_OP_1001J1_64_4995_n422 ) 
    , .CO ( DP_OP_1001J1_64_4995_n406 ) , .S ( DP_OP_1001J1_64_4995_n407 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U302 (.A ( in_reg_salida_v[5] ) 
    , .B ( coeficiente_a22_in[11] ) , .CI ( coeficiente_a22_in[9] ) 
    , .CO ( DP_OP_1001J1_64_4995_n424 ) , .S ( DP_OP_1001J1_64_4995_n425 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U326 (.A ( DP_OP_1001J1_64_4995_n482 ) 
    , .B ( DP_OP_1001J1_64_4995_n480 ) , .CI ( DP_OP_1001J1_64_4995_n479 ) 
    , .CO ( DP_OP_1001J1_64_4995_n470 ) , .S ( DP_OP_1001J1_64_4995_n471 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U273 (.A ( n1587 ) , .B ( n1533 ) 
    , .CI ( sos2_reg_entrada[18] ) , .CO ( DP_OP_1001J1_64_4995_n366 ) 
    , .S ( DP_OP_1001J1_64_4995_n367 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U295 (.A ( sos2_reg_entrada[14] ) 
    , .B ( in_reg_salida_v[6] ) , .CI ( coeficiente_a22_in[12] ) 
    , .CO ( DP_OP_1001J1_64_4995_n410 ) , .S ( DP_OP_1001J1_64_4995_n411 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U149 (.A ( n1553 ) 
    , .B ( DP_OP_1001J1_64_4995_n274 ) , .CI ( DP_OP_1001J1_64_4995_n550 ) 
    , .CO ( DP_OP_1001J1_64_4995_n187 ) , .S ( partial_2_L[0] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U255 (.A ( DP_OP_1001J1_64_4995_n485 ) 
    , .B ( DP_OP_1001J1_64_4995_n483 ) , .CI ( DP_OP_1001J1_64_4995_n481 ) 
    , .CO ( DP_OP_1001J1_64_4995_n333 ) , .S ( partial_1[0] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U318 (.A ( DP_OP_1001J1_64_4995_n463 ) 
    , .B ( DP_OP_1001J1_64_4995_n472 ) , .CI ( DP_OP_1001J1_64_4995_n470 ) 
    , .CO ( DP_OP_1001J1_64_4995_n456 ) , .S ( DP_OP_1001J1_64_4995_n457 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U171 (.A ( coeficiente_b12_L_v_out[9] ) 
    , .B ( n1557 ) , .CI ( coeficiente_b11_L_v_out[18] ) 
    , .CO ( DP_OP_1001J1_64_4995_n227 ) , .S ( DP_OP_1001J1_64_4995_n228 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U328 (.A ( n1585 ) , .B ( n1584 ) , .CI ( n1542 ) 
    , .CO ( DP_OP_1001J1_64_4995_n474 ) , .S ( DP_OP_1001J1_64_4995_n475 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U321 (.A ( n1581 ) , .B ( n1584 ) , .CI ( n1543 ) 
    , .CO ( DP_OP_1001J1_64_4995_n462 ) , .S ( DP_OP_1001J1_64_4995_n463 ) ) ;
HADDX1 DP_OP_1001J1_64_4995_U330 (.B0 ( in_reg_salida_v[1] ) 
    , .A0 ( coeficiente_a22_in[5] ) , .C1 ( DP_OP_1001J1_64_4995_n478 ) 
    , .SO ( DP_OP_1001J1_64_4995_n479 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U301 (.A ( n1546 ) , .B ( n1560 ) , .CI ( n1584 ) 
    , .CO ( DP_OP_1001J1_64_4995_n422 ) , .S ( DP_OP_1001J1_64_4995_n423 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U288 (.A ( in_reg_salida_v[7] ) , .B ( n1548 ) 
    , .CI ( n1585 ) , .CO ( DP_OP_1001J1_64_4995_n396 ) 
    , .S ( DP_OP_1001J1_64_4995_n397 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U315 (.A ( coeficiente_a22_in[9] ) , .B ( n1560 ) 
    , .CI ( n1582 ) , .CO ( DP_OP_1001J1_64_4995_n450 ) 
    , .S ( DP_OP_1001J1_64_4995_n451 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U308 (.A ( coeficiente_a22_in[10] ) , .B ( n1587 ) 
    , .CI ( n1583 ) , .CO ( DP_OP_1001J1_64_4995_n436 ) 
    , .S ( DP_OP_1001J1_64_4995_n437 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U162 (.A ( coeficiente_b12_L_v_out[12] ) 
    , .B ( n1513 ) , .CI ( DP_OP_1001J1_64_4995_n213 ) 
    , .CO ( DP_OP_1001J1_64_4995_n209 ) , .S ( DP_OP_1001J1_64_4995_n210 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U168 (.A ( n1507 ) 
    , .B ( DP_OP_1001J1_64_4995_n227 ) , .CI ( DP_OP_1001J1_64_4995_n225 ) 
    , .CO ( DP_OP_1001J1_64_4995_n221 ) , .S ( DP_OP_1001J1_64_4995_n222 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U170 (.A ( DP_OP_1001J1_64_4995_n228 ) 
    , .B ( DP_OP_1001J1_64_4995_n231 ) , .CI ( DP_OP_1001J1_64_4995_n229 ) 
    , .CO ( DP_OP_1001J1_64_4995_n225 ) , .S ( DP_OP_1001J1_64_4995_n226 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U172 (.A ( DP_OP_1001J1_64_4995_n235 ) 
    , .B ( DP_OP_1001J1_64_4995_n232 ) , .CI ( DP_OP_1001J1_64_4995_n233 ) 
    , .CO ( DP_OP_1001J1_64_4995_n229 ) , .S ( DP_OP_1001J1_64_4995_n230 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U174 (.A ( DP_OP_1001J1_64_4995_n241 ) 
    , .B ( DP_OP_1001J1_64_4995_n236 ) , .CI ( DP_OP_1001J1_64_4995_n239 ) 
    , .CO ( DP_OP_1001J1_64_4995_n233 ) , .S ( DP_OP_1001J1_64_4995_n234 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U177 (.A ( DP_OP_1001J1_64_4995_n247 ) 
    , .B ( DP_OP_1001J1_64_4995_n242 ) , .CI ( DP_OP_1001J1_64_4995_n245 ) 
    , .CO ( DP_OP_1001J1_64_4995_n239 ) , .S ( DP_OP_1001J1_64_4995_n240 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U180 (.A ( DP_OP_1001J1_64_4995_n253 ) 
    , .B ( DP_OP_1001J1_64_4995_n248 ) , .CI ( DP_OP_1001J1_64_4995_n251 ) 
    , .CO ( DP_OP_1001J1_64_4995_n245 ) , .S ( DP_OP_1001J1_64_4995_n246 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U175 (.A ( n1558 ) 
    , .B ( DP_OP_1001J1_64_4995_n243 ) , .CI ( DP_OP_1001J1_64_4995_n238 ) 
    , .CO ( DP_OP_1001J1_64_4995_n235 ) , .S ( DP_OP_1001J1_64_4995_n236 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U176 (.A ( coeficiente_b12_L_v_out[7] ) 
    , .B ( n1555 ) , .CI ( n1556 ) , .CO ( DP_OP_1001J1_64_4995_n237 ) 
    , .S ( DP_OP_1001J1_64_4995_n238 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U178 (.A ( n1554 ) 
    , .B ( DP_OP_1001J1_64_4995_n249 ) , .CI ( DP_OP_1001J1_64_4995_n244 ) 
    , .CO ( DP_OP_1001J1_64_4995_n241 ) , .S ( DP_OP_1001J1_64_4995_n242 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U183 (.A ( DP_OP_1001J1_64_4995_n259 ) 
    , .B ( DP_OP_1001J1_64_4995_n254 ) , .CI ( DP_OP_1001J1_64_4995_n257 ) 
    , .CO ( DP_OP_1001J1_64_4995_n251 ) , .S ( DP_OP_1001J1_64_4995_n252 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U184 (.A ( n1557 ) 
    , .B ( DP_OP_1001J1_64_4995_n261 ) , .CI ( DP_OP_1001J1_64_4995_n256 ) 
    , .CO ( DP_OP_1001J1_64_4995_n253 ) , .S ( DP_OP_1001J1_64_4995_n254 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U154 (.A ( coeficiente_b12_L_v_out[16] ) 
    , .B ( n1521 ) , .CI ( DP_OP_1001J1_64_4995_n197 ) 
    , .CO ( DP_OP_1001J1_64_4995_n193 ) , .S ( DP_OP_1001J1_64_4995_n194 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U156 (.A ( coeficiente_b12_L_v_out[15] ) 
    , .B ( n1519 ) , .CI ( DP_OP_1001J1_64_4995_n201 ) 
    , .CO ( DP_OP_1001J1_64_4995_n197 ) , .S ( DP_OP_1001J1_64_4995_n198 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U158 (.A ( coeficiente_b12_L_v_out[14] ) 
    , .B ( n1517 ) , .CI ( DP_OP_1001J1_64_4995_n205 ) 
    , .CO ( DP_OP_1001J1_64_4995_n201 ) , .S ( DP_OP_1001J1_64_4995_n202 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U160 (.A ( coeficiente_b12_L_v_out[13] ) 
    , .B ( n1515 ) , .CI ( DP_OP_1001J1_64_4995_n209 ) 
    , .CO ( DP_OP_1001J1_64_4995_n205 ) , .S ( DP_OP_1001J1_64_4995_n206 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U73 (.A ( DP_OP_1001J1_64_4995_n106 ) 
    , .B ( DP_OP_1001J1_64_4995_n101 ) , .CI ( DP_OP_1001J1_64_4995_n104 ) 
    , .CO ( DP_OP_1001J1_64_4995_n98 ) , .S ( DP_OP_1001J1_64_4995_n99 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U194 (.A ( coeficiente_b12_L_v_out[0] ) 
    , .B ( coeficiente_b11_L_v_out[11] ) , .CI ( n1559 ) 
    , .CO ( DP_OP_1001J1_64_4995_n273 ) , .S ( DP_OP_1001J1_64_4995_n274 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U193 (.A ( coeficiente_b12_L_v_out[1] ) 
    , .B ( coeficiente_b11_L_v_out[10] ) , .CI ( coeficiente_b11_L_v_out[12] ) 
    , .CO ( DP_OP_1001J1_64_4995_n271 ) , .S ( DP_OP_1001J1_64_4995_n272 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U191 (.A ( coeficiente_b12_L_v_out[2] ) 
    , .B ( coeficiente_b11_L_v_out[13] ) , .CI ( n1551 ) 
    , .CO ( DP_OP_1001J1_64_4995_n267 ) , .S ( DP_OP_1001J1_64_4995_n268 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U189 (.A ( DP_OP_1001J1_64_4995_n268 ) 
    , .B ( DP_OP_1001J1_64_4995_n269 ) , .CI ( DP_OP_1001J1_64_4995_n266 ) 
    , .CO ( DP_OP_1001J1_64_4995_n263 ) , .S ( DP_OP_1001J1_64_4995_n264 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U190 (.A ( n1555 ) , .B ( n1550 ) 
    , .CI ( DP_OP_1001J1_64_4995_n271 ) , .CO ( DP_OP_1001J1_64_4995_n265 ) 
    , .S ( DP_OP_1001J1_64_4995_n266 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U186 (.A ( DP_OP_1001J1_64_4995_n265 ) 
    , .B ( DP_OP_1001J1_64_4995_n260 ) , .CI ( DP_OP_1001J1_64_4995_n263 ) 
    , .CO ( DP_OP_1001J1_64_4995_n257 ) , .S ( DP_OP_1001J1_64_4995_n258 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U187 (.A ( n1556 ) 
    , .B ( DP_OP_1001J1_64_4995_n267 ) , .CI ( DP_OP_1001J1_64_4995_n262 ) 
    , .CO ( DP_OP_1001J1_64_4995_n259 ) , .S ( DP_OP_1001J1_64_4995_n260 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U79 (.A ( DP_OP_1001J1_64_4995_n118 ) 
    , .B ( DP_OP_1001J1_64_4995_n113 ) , .CI ( DP_OP_1001J1_64_4995_n116 ) 
    , .CO ( DP_OP_1001J1_64_4995_n110 ) , .S ( DP_OP_1001J1_64_4995_n111 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U66 (.A ( coeficiente_b12_H_v_out[8] ) 
    , .B ( coeficiente_a11_H_in[17] ) , .CI ( DP_OP_1001J1_64_4995_n90 ) 
    , .CO ( DP_OP_1001J1_64_4995_n84 ) , .S ( DP_OP_1001J1_64_4995_n85 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U76 (.A ( DP_OP_1001J1_64_4995_n112 ) 
    , .B ( DP_OP_1001J1_64_4995_n107 ) , .CI ( DP_OP_1001J1_64_4995_n110 ) 
    , .CO ( DP_OP_1001J1_64_4995_n104 ) , .S ( DP_OP_1001J1_64_4995_n105 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U61 (.A ( n1508 ) 
    , .B ( DP_OP_1001J1_64_4995_n80 ) , .CI ( DP_OP_1001J1_64_4995_n78 ) 
    , .CO ( DP_OP_1001J1_64_4995_n74 ) , .S ( DP_OP_1001J1_64_4995_n75 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U63 (.A ( DP_OP_1001J1_64_4995_n81 ) 
    , .B ( DP_OP_1001J1_64_4995_n84 ) , .CI ( DP_OP_1001J1_64_4995_n82 ) 
    , .CO ( DP_OP_1001J1_64_4995_n78 ) , .S ( DP_OP_1001J1_64_4995_n79 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U65 (.A ( DP_OP_1001J1_64_4995_n88 ) 
    , .B ( DP_OP_1001J1_64_4995_n85 ) , .CI ( DP_OP_1001J1_64_4995_n86 ) 
    , .CO ( DP_OP_1001J1_64_4995_n82 ) , .S ( DP_OP_1001J1_64_4995_n83 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U67 (.A ( DP_OP_1001J1_64_4995_n94 ) 
    , .B ( DP_OP_1001J1_64_4995_n89 ) , .CI ( DP_OP_1001J1_64_4995_n92 ) 
    , .CO ( DP_OP_1001J1_64_4995_n86 ) , .S ( DP_OP_1001J1_64_4995_n87 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U70 (.A ( DP_OP_1001J1_64_4995_n100 ) 
    , .B ( DP_OP_1001J1_64_4995_n95 ) , .CI ( DP_OP_1001J1_64_4995_n98 ) 
    , .CO ( DP_OP_1001J1_64_4995_n92 ) , .S ( DP_OP_1001J1_64_4995_n93 ) ) ;
DFFNX1 secuencia_reloj_prioridad_salida_reg_0_ (
    .CLK ( filtro_pipelining_clk_2x ) 
    , .D ( secuencia_reloj_prioridad_salida_pre_0_ ) , .QN ( n1035 ) 
    , .Q ( n1492 ) ) ;
DFFNX1 secuencia_reloj_prioridad_salida_reg_2_ (
    .CLK ( filtro_pipelining_clk_2x ) , .D ( n1120 ) , .QN ( seleccion_2_ ) 
    , .Q ( n1493 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U87 (.A ( coeficiente_b12_H_v_out[0] ) 
    , .B ( coeficiente_a11_H_in[11] ) , .CI ( n1502 ) 
    , .CO ( DP_OP_1001J1_64_4995_n126 ) , .S ( DP_OP_1001J1_64_4995_n127 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U86 (.A ( coeficiente_b12_H_v_out[1] ) 
    , .B ( coeficiente_a11_H_in[10] ) , .CI ( coeficiente_a11_H_in[12] ) 
    , .CO ( DP_OP_1001J1_64_4995_n124 ) , .S ( DP_OP_1001J1_64_4995_n125 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U84 (.A ( coeficiente_b12_H_v_out[2] ) 
    , .B ( coeficiente_a11_H_in[13] ) , .CI ( n1524 ) 
    , .CO ( DP_OP_1001J1_64_4995_n120 ) , .S ( DP_OP_1001J1_64_4995_n121 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U81 (.A ( coeficiente_b12_H_v_out[3] ) 
    , .B ( coeficiente_a11_H_in[14] ) , .CI ( n1525 ) 
    , .CO ( DP_OP_1001J1_64_4995_n114 ) , .S ( DP_OP_1001J1_64_4995_n115 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U78 (.A ( coeficiente_b12_H_v_out[4] ) 
    , .B ( coeficiente_a11_H_in[15] ) , .CI ( n1526 ) 
    , .CO ( DP_OP_1001J1_64_4995_n108 ) , .S ( DP_OP_1001J1_64_4995_n109 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U82 (.A ( DP_OP_1001J1_64_4995_n121 ) 
    , .B ( DP_OP_1001J1_64_4995_n122 ) , .CI ( DP_OP_1001J1_64_4995_n119 ) 
    , .CO ( DP_OP_1001J1_64_4995_n116 ) , .S ( DP_OP_1001J1_64_4995_n117 ) ) ;
INVX0 U6 (.ZN ( n1034 ) , .INP ( reloj_secuencia[5] ) ) ;
DFFNX1 reloj_secuencia_delay_reg_0_ (.CLK ( filtro_pipelining_clk_2x ) 
    , .D ( reloj_secuencia[0] ) , .Q ( reloj_secuencia_delay[0] ) ) ;
DFFNX1 reloj_secuencia_delay_reg_1_ (.CLK ( filtro_pipelining_clk_2x ) 
    , .D ( reloj_secuencia[1] ) , .Q ( reloj_secuencia_delay[1] ) ) ;
DFFNX1 reloj_secuencia_delay_reg_2_ (.CLK ( filtro_pipelining_clk_2x ) 
    , .D ( reloj_secuencia[2] ) , .Q ( reloj_secuencia_delay[2] ) ) ;
DFFNX1 reloj_secuencia_delay_reg_3_ (.CLK ( filtro_pipelining_clk_2x ) 
    , .D ( reloj_secuencia[3] ) , .Q ( reloj_secuencia_delay[3] ) ) ;
DFFNX1 reloj_secuencia_delay_reg_4_ (.CLK ( filtro_pipelining_clk_2x ) 
    , .D ( reloj_secuencia[4] ) , .Q ( reloj_secuencia_delay[4] ) ) ;
DFFNX1 reloj_secuencia_delay_reg_6_ (.CLK ( filtro_pipelining_clk_2x ) 
    , .D ( reloj_secuencia[6] ) , .Q ( reloj_secuencia_delay[6] ) ) ;
DFFNX1 reloj_secuencia_delay_reg_5_ (.CLK ( filtro_pipelining_clk_2x ) 
    , .D ( n1034 ) , .QN ( reloj_secuencia_delay[5] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U136 (.A ( DP_OP_1001J1_64_4995_n210 ) 
    , .B ( DP_OP_1001J1_64_4995_n563 ) , .CI ( DP_OP_1001J1_64_4995_n175 ) 
    , .CO ( DP_OP_1001J1_64_4995_n174 ) , .S ( partial_2_L[13] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U137 (.A ( DP_OP_1001J1_64_4995_n214 ) 
    , .B ( DP_OP_1001J1_64_4995_n562 ) , .CI ( DP_OP_1001J1_64_4995_n176 ) 
    , .CO ( DP_OP_1001J1_64_4995_n175 ) , .S ( partial_2_L[12] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U239 (.A ( DP_OP_1001J1_64_4995_n339 ) 
    , .B ( DP_OP_1001J1_64_4995_n340 ) , .CI ( DP_OP_1001J1_64_4995_n318 ) 
    , .CO ( DP_OP_1001J1_64_4995_n317 ) , .S ( partial_1[16] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U242 (.A ( DP_OP_1001J1_64_4995_n350 ) 
    , .B ( DP_OP_1001J1_64_4995_n347 ) , .CI ( DP_OP_1001J1_64_4995_n321 ) 
    , .CO ( DP_OP_1001J1_64_4995_n320 ) , .S ( partial_1[13] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U243 (.A ( DP_OP_1001J1_64_4995_n356 ) 
    , .B ( DP_OP_1001J1_64_4995_n351 ) , .CI ( DP_OP_1001J1_64_4995_n322 ) 
    , .CO ( DP_OP_1001J1_64_4995_n321 ) , .S ( partial_1[12] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U244 (.A ( DP_OP_1001J1_64_4995_n357 ) 
    , .B ( DP_OP_1001J1_64_4995_n362 ) , .CI ( DP_OP_1001J1_64_4995_n323 ) 
    , .CO ( DP_OP_1001J1_64_4995_n322 ) , .S ( partial_1[11] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U245 (.A ( DP_OP_1001J1_64_4995_n370 ) 
    , .B ( DP_OP_1001J1_64_4995_n363 ) , .CI ( DP_OP_1001J1_64_4995_n324 ) 
    , .CO ( DP_OP_1001J1_64_4995_n323 ) , .S ( partial_1[10] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U238 (.A ( DP_OP_1001J1_64_4995_n338 ) 
    , .B ( DP_OP_1001J1_64_4995_n337 ) , .CI ( DP_OP_1001J1_64_4995_n317 ) 
    , .CO ( DP_OP_1001J1_64_4995_n316 ) , .S ( partial_1[17] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U26 (.A ( DP_OP_1001J1_64_4995_n51 ) 
    , .B ( DP_OP_1001J1_64_4995_n566 ) , .CI ( DP_OP_1001J1_64_4995_n25 ) 
    , .CO ( DP_OP_1001J1_64_4995_n24 ) , .S ( partial_2_H[16] ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U6 (.A ( DP_OP_1003J1_66_5789_n24 ) 
    , .B ( DP_OP_1003J1_66_5789_n25 ) , .CI ( DP_OP_1003J1_66_5789_n6 ) 
    , .CO ( DP_OP_1003J1_66_5789_n5 ) , .S ( bajo_reg_entrada[13] ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U7 (.A ( DP_OP_1003J1_66_5789_n27 ) 
    , .B ( DP_OP_1003J1_66_5789_n26 ) , .CI ( DP_OP_1003J1_66_5789_n7 ) 
    , .CO ( DP_OP_1003J1_66_5789_n6 ) , .S ( bajo_reg_entrada[12] ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U8 (.A ( DP_OP_1003J1_66_5789_n31 ) 
    , .B ( DP_OP_1003J1_66_5789_n28 ) , .CI ( DP_OP_1003J1_66_5789_n8 ) 
    , .CO ( DP_OP_1003J1_66_5789_n7 ) , .S ( bajo_reg_entrada[11] ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U9 (.A ( DP_OP_1003J1_66_5789_n35 ) 
    , .B ( DP_OP_1003J1_66_5789_n32 ) , .CI ( DP_OP_1003J1_66_5789_n9 ) 
    , .CO ( DP_OP_1003J1_66_5789_n8 ) , .S ( bajo_reg_entrada[10] ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U10 (.A ( DP_OP_1003J1_66_5789_n39 ) 
    , .B ( DP_OP_1003J1_66_5789_n36 ) , .CI ( DP_OP_1003J1_66_5789_n10 ) 
    , .CO ( DP_OP_1003J1_66_5789_n9 ) , .S ( bajo_reg_entrada[9] ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U11 (.A ( DP_OP_1003J1_66_5789_n43 ) 
    , .B ( DP_OP_1003J1_66_5789_n40 ) , .CI ( DP_OP_1003J1_66_5789_n11 ) 
    , .CO ( DP_OP_1003J1_66_5789_n10 ) , .S ( bajo_reg_entrada[8] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U132 (.A ( DP_OP_1001J1_64_4995_n194 ) 
    , .B ( DP_OP_1001J1_64_4995_n567 ) , .CI ( DP_OP_1001J1_64_4995_n171 ) 
    , .CO ( DP_OP_1001J1_64_4995_n170 ) , .S ( partial_2_L[17] ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U6 (.A ( DP_OP_1004J1_67_3033_n24 ) 
    , .B ( DP_OP_1004J1_67_3033_n25 ) , .CI ( DP_OP_1004J1_67_3033_n6 ) 
    , .CO ( DP_OP_1004J1_67_3033_n5 ) , .S ( alto_reg_entrada[13] ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U7 (.A ( DP_OP_1004J1_67_3033_n27 ) 
    , .B ( DP_OP_1004J1_67_3033_n26 ) , .CI ( DP_OP_1004J1_67_3033_n7 ) 
    , .CO ( DP_OP_1004J1_67_3033_n6 ) , .S ( alto_reg_entrada[12] ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U8 (.A ( DP_OP_1004J1_67_3033_n31 ) 
    , .B ( DP_OP_1004J1_67_3033_n28 ) , .CI ( DP_OP_1004J1_67_3033_n8 ) 
    , .CO ( DP_OP_1004J1_67_3033_n7 ) , .S ( alto_reg_entrada[11] ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U10 (.A ( DP_OP_1004J1_67_3033_n39 ) 
    , .B ( DP_OP_1004J1_67_3033_n36 ) , .CI ( DP_OP_1004J1_67_3033_n10 ) 
    , .CO ( DP_OP_1004J1_67_3033_n9 ) , .S ( alto_reg_entrada[9] ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U18 (.A ( DP_OP_1004J1_67_3033_n82 ) 
    , .B ( DP_OP_1004J1_67_3033_n18 ) , .CI ( DP_OP_1004J1_67_3033_n80 ) 
    , .CO ( DP_OP_1004J1_67_3033_n17 ) , .S ( alto_reg_entrada[1] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U4 (.A ( coeficiente_b11_H_v_out[17] ) 
    , .B ( partial_2_H[17] ) , .CI ( DP_OP_1001J1_64_4995_n4 ) 
    , .CO ( DP_OP_1001J1_64_4995_n3 ) , .S ( partial_3_H[17] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U25 (.A ( DP_OP_1001J1_64_4995_n47 ) 
    , .B ( DP_OP_1001J1_64_4995_n567 ) , .CI ( DP_OP_1001J1_64_4995_n24 ) 
    , .CO ( DP_OP_1001J1_64_4995_n23 ) , .S ( partial_2_H[17] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U5 (.A ( coeficiente_b11_H_v_out[16] ) 
    , .B ( partial_2_H[16] ) , .CI ( DP_OP_1001J1_64_4995_n5 ) 
    , .CO ( DP_OP_1001J1_64_4995_n4 ) , .S ( partial_3_H[16] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U41 (.A ( DP_OP_1001J1_64_4995_n123 ) 
    , .B ( DP_OP_1001J1_64_4995_n40 ) , .CI ( DP_OP_1001J1_64_4995_n551 ) 
    , .CO ( DP_OP_1001J1_64_4995_n39 ) , .S ( partial_2_H[1] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U148 (.A ( DP_OP_1001J1_64_4995_n270 ) 
    , .B ( DP_OP_1001J1_64_4995_n187 ) , .CI ( DP_OP_1001J1_64_4995_n551 ) 
    , .CO ( DP_OP_1001J1_64_4995_n186 ) , .S ( partial_2_L[1] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U252 (.A ( DP_OP_1001J1_64_4995_n454 ) 
    , .B ( DP_OP_1001J1_64_4995_n441 ) , .CI ( DP_OP_1001J1_64_4995_n331 ) 
    , .CO ( DP_OP_1001J1_64_4995_n330 ) , .S ( partial_1[3] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U253 (.A ( DP_OP_1001J1_64_4995_n457 ) 
    , .B ( DP_OP_1001J1_64_4995_n455 ) , .CI ( DP_OP_1001J1_64_4995_n332 ) 
    , .CO ( DP_OP_1001J1_64_4995_n331 ) , .S ( partial_1[2] ) ) ;
HADDX1 DP_OP_1001J1_64_4995_U235 (.B0 ( coeficiente_a22_in[0] ) 
    , .A0 ( partial_1[0] ) , .C1 ( DP_OP_1001J1_64_4995_n314 ) 
    , .SO ( DP_OP_1001J1_64_4995_n550 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U254 (.A ( DP_OP_1001J1_64_4995_n333 ) 
    , .B ( DP_OP_1001J1_64_4995_n471 ) , .CI ( DP_OP_1001J1_64_4995_n469 ) 
    , .CO ( DP_OP_1001J1_64_4995_n332 ) , .S ( partial_1[1] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U332 (.A ( sos2_reg_entrada[13] ) 
    , .B ( in_reg_salida_v[0] ) , .CI ( n1541 ) 
    , .CO ( DP_OP_1001J1_64_4995_n482 ) , .S ( DP_OP_1001J1_64_4995_n483 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U333 (.A ( coeficiente_a22_in[13] ) 
    , .B ( coeficiente_a22_in[6] ) , .CI ( coeficiente_a22_in[4] ) 
    , .CO ( DP_OP_1001J1_64_4995_n484 ) , .S ( DP_OP_1001J1_64_4995_n485 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U226 (.A ( coeficiente_a22_in[9] ) 
    , .B ( partial_1[9] ) , .CI ( DP_OP_1001J1_64_4995_n306 ) 
    , .CO ( DP_OP_1001J1_64_4995_n305 ) , .S ( DP_OP_1001J1_64_4995_n559 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U227 (.A ( coeficiente_a22_in[8] ) 
    , .B ( partial_1[8] ) , .CI ( DP_OP_1001J1_64_4995_n307 ) 
    , .CO ( DP_OP_1001J1_64_4995_n306 ) , .S ( DP_OP_1001J1_64_4995_n558 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U246 (.A ( DP_OP_1001J1_64_4995_n378 ) 
    , .B ( DP_OP_1001J1_64_4995_n371 ) , .CI ( DP_OP_1001J1_64_4995_n325 ) 
    , .CO ( DP_OP_1001J1_64_4995_n324 ) , .S ( partial_1[9] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U39 (.A ( DP_OP_1001J1_64_4995_n111 ) 
    , .B ( DP_OP_1001J1_64_4995_n38 ) , .CI ( DP_OP_1001J1_64_4995_n553 ) 
    , .CO ( DP_OP_1001J1_64_4995_n37 ) , .S ( partial_2_H[3] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U247 (.A ( DP_OP_1001J1_64_4995_n388 ) 
    , .B ( DP_OP_1001J1_64_4995_n379 ) , .CI ( DP_OP_1001J1_64_4995_n326 ) 
    , .CO ( DP_OP_1001J1_64_4995_n325 ) , .S ( partial_1[8] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U146 (.A ( DP_OP_1001J1_64_4995_n258 ) 
    , .B ( DP_OP_1001J1_64_4995_n185 ) , .CI ( DP_OP_1001J1_64_4995_n553 ) 
    , .CO ( DP_OP_1001J1_64_4995_n184 ) , .S ( partial_2_L[3] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U40 (.A ( DP_OP_1001J1_64_4995_n117 ) 
    , .B ( DP_OP_1001J1_64_4995_n39 ) , .CI ( DP_OP_1001J1_64_4995_n552 ) 
    , .CO ( DP_OP_1001J1_64_4995_n38 ) , .S ( partial_2_H[2] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U147 (.A ( DP_OP_1001J1_64_4995_n264 ) 
    , .B ( DP_OP_1001J1_64_4995_n186 ) , .CI ( DP_OP_1001J1_64_4995_n552 ) 
    , .CO ( DP_OP_1001J1_64_4995_n185 ) , .S ( partial_2_L[2] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U33 (.A ( DP_OP_1001J1_64_4995_n79 ) 
    , .B ( DP_OP_1001J1_64_4995_n559 ) , .CI ( DP_OP_1001J1_64_4995_n32 ) 
    , .CO ( DP_OP_1001J1_64_4995_n31 ) , .S ( partial_2_H[9] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U139 (.A ( DP_OP_1001J1_64_4995_n222 ) 
    , .B ( DP_OP_1001J1_64_4995_n560 ) , .CI ( DP_OP_1001J1_64_4995_n178 ) 
    , .CO ( DP_OP_1001J1_64_4995_n177 ) , .S ( partial_2_L[10] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U222 (.A ( coeficiente_a22_in[13] ) 
    , .B ( partial_1[13] ) , .CI ( DP_OP_1001J1_64_4995_n302 ) 
    , .CO ( DP_OP_1001J1_64_4995_n301 ) , .S ( DP_OP_1001J1_64_4995_n563 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U140 (.A ( DP_OP_1001J1_64_4995_n226 ) 
    , .B ( DP_OP_1001J1_64_4995_n559 ) , .CI ( DP_OP_1001J1_64_4995_n179 ) 
    , .CO ( DP_OP_1001J1_64_4995_n178 ) , .S ( partial_2_L[9] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U223 (.A ( coeficiente_a22_in[12] ) 
    , .B ( partial_1[12] ) , .CI ( DP_OP_1001J1_64_4995_n303 ) 
    , .CO ( DP_OP_1001J1_64_4995_n302 ) , .S ( DP_OP_1001J1_64_4995_n562 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U224 (.A ( coeficiente_a22_in[11] ) 
    , .B ( partial_1[11] ) , .CI ( DP_OP_1001J1_64_4995_n304 ) 
    , .CO ( DP_OP_1001J1_64_4995_n303 ) , .S ( DP_OP_1001J1_64_4995_n561 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U141 (.A ( DP_OP_1001J1_64_4995_n230 ) 
    , .B ( DP_OP_1001J1_64_4995_n558 ) , .CI ( DP_OP_1001J1_64_4995_n180 ) 
    , .CO ( DP_OP_1001J1_64_4995_n179 ) , .S ( partial_2_L[8] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U225 (.A ( coeficiente_a22_in[10] ) 
    , .B ( partial_1[10] ) , .CI ( DP_OP_1001J1_64_4995_n305 ) 
    , .CO ( DP_OP_1001J1_64_4995_n304 ) , .S ( DP_OP_1001J1_64_4995_n560 ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U29 (.A ( DP_OP_1001J1_64_4995_n63 ) 
    , .B ( DP_OP_1001J1_64_4995_n563 ) , .CI ( DP_OP_1001J1_64_4995_n28 ) 
    , .CO ( DP_OP_1001J1_64_4995_n27 ) , .S ( partial_2_H[13] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U30 (.A ( DP_OP_1001J1_64_4995_n67 ) 
    , .B ( DP_OP_1001J1_64_4995_n562 ) , .CI ( DP_OP_1001J1_64_4995_n29 ) 
    , .CO ( DP_OP_1001J1_64_4995_n28 ) , .S ( partial_2_H[12] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U117 (.A ( coeficiente_b11_L_v_out[11] ) 
    , .B ( partial_2_L[11] ) , .CI ( DP_OP_1001J1_64_4995_n157 ) 
    , .CO ( DP_OP_1001J1_64_4995_n156 ) , .S ( partial_3_L[11] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U31 (.A ( DP_OP_1001J1_64_4995_n71 ) 
    , .B ( DP_OP_1001J1_64_4995_n561 ) , .CI ( DP_OP_1001J1_64_4995_n30 ) 
    , .CO ( DP_OP_1001J1_64_4995_n29 ) , .S ( partial_2_H[11] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U240 (.A ( DP_OP_1001J1_64_4995_n342 ) 
    , .B ( DP_OP_1001J1_64_4995_n341 ) , .CI ( DP_OP_1001J1_64_4995_n319 ) 
    , .CO ( DP_OP_1001J1_64_4995_n318 ) , .S ( partial_1[15] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U118 (.A ( coeficiente_b11_L_v_out[10] ) 
    , .B ( partial_2_L[10] ) , .CI ( DP_OP_1001J1_64_4995_n158 ) 
    , .CO ( DP_OP_1001J1_64_4995_n157 ) , .S ( partial_3_L[10] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U138 (.A ( DP_OP_1001J1_64_4995_n218 ) 
    , .B ( DP_OP_1001J1_64_4995_n561 ) , .CI ( DP_OP_1001J1_64_4995_n177 ) 
    , .CO ( DP_OP_1001J1_64_4995_n176 ) , .S ( partial_2_L[11] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U241 (.A ( DP_OP_1001J1_64_4995_n346 ) 
    , .B ( DP_OP_1001J1_64_4995_n343 ) , .CI ( DP_OP_1001J1_64_4995_n320 ) 
    , .CO ( DP_OP_1001J1_64_4995_n319 ) , .S ( partial_1[14] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U133 (.A ( DP_OP_1001J1_64_4995_n198 ) 
    , .B ( DP_OP_1001J1_64_4995_n566 ) , .CI ( DP_OP_1001J1_64_4995_n172 ) 
    , .CO ( DP_OP_1001J1_64_4995_n171 ) , .S ( partial_2_L[16] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U27 (.A ( DP_OP_1001J1_64_4995_n55 ) 
    , .B ( DP_OP_1001J1_64_4995_n565 ) , .CI ( DP_OP_1001J1_64_4995_n26 ) 
    , .CO ( DP_OP_1001J1_64_4995_n25 ) , .S ( partial_2_H[15] ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U17 (.A ( DP_OP_1003J1_66_5789_n67 ) 
    , .B ( DP_OP_1003J1_66_5789_n64 ) , .CI ( DP_OP_1003J1_66_5789_n17 ) 
    , .CO ( DP_OP_1003J1_66_5789_n16 ) , .S ( bajo_reg_entrada[2] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U8 (.A ( coeficiente_b11_H_v_out[13] ) 
    , .B ( partial_2_H[13] ) , .CI ( DP_OP_1001J1_64_4995_n8 ) 
    , .CO ( DP_OP_1001J1_64_4995_n7 ) , .S ( partial_3_H[13] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U28 (.A ( DP_OP_1001J1_64_4995_n59 ) 
    , .B ( DP_OP_1001J1_64_4995_n564 ) , .CI ( DP_OP_1001J1_64_4995_n27 ) 
    , .CO ( DP_OP_1001J1_64_4995_n26 ) , .S ( partial_2_H[14] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U134 (.A ( DP_OP_1001J1_64_4995_n202 ) 
    , .B ( DP_OP_1001J1_64_4995_n565 ) , .CI ( DP_OP_1001J1_64_4995_n173 ) 
    , .CO ( DP_OP_1001J1_64_4995_n172 ) , .S ( partial_2_L[15] ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U18 (.A ( DP_OP_1003J1_66_5789_n70 ) 
    , .B ( DP_OP_1003J1_66_5789_n18 ) , .CI ( DP_OP_1003J1_66_5789_n68 ) 
    , .CO ( DP_OP_1003J1_66_5789_n17 ) , .S ( bajo_reg_entrada[1] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U135 (.A ( DP_OP_1001J1_64_4995_n206 ) 
    , .B ( DP_OP_1001J1_64_4995_n564 ) , .CI ( DP_OP_1001J1_64_4995_n174 ) 
    , .CO ( DP_OP_1001J1_64_4995_n173 ) , .S ( partial_2_L[14] ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U9 (.A ( DP_OP_1004J1_67_3033_n35 ) 
    , .B ( DP_OP_1004J1_67_3033_n32 ) , .CI ( DP_OP_1004J1_67_3033_n9 ) 
    , .CO ( DP_OP_1004J1_67_3033_n8 ) , .S ( alto_reg_entrada[10] ) ) ;
FADDX1 DP_OP_1004J1_67_3033_U17 (.A ( DP_OP_1004J1_67_3033_n79 ) 
    , .B ( DP_OP_1004J1_67_3033_n74 ) , .CI ( DP_OP_1004J1_67_3033_n17 ) 
    , .CO ( DP_OP_1004J1_67_3033_n16 ) , .S ( alto_reg_entrada[2] ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U12 (.A ( DP_OP_1003J1_66_5789_n47 ) 
    , .B ( DP_OP_1003J1_66_5789_n44 ) , .CI ( DP_OP_1003J1_66_5789_n12 ) 
    , .CO ( DP_OP_1003J1_66_5789_n11 ) , .S ( bajo_reg_entrada[7] ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U13 (.A ( DP_OP_1003J1_66_5789_n51 ) 
    , .B ( DP_OP_1003J1_66_5789_n48 ) , .CI ( DP_OP_1003J1_66_5789_n13 ) 
    , .CO ( DP_OP_1003J1_66_5789_n12 ) , .S ( bajo_reg_entrada[6] ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U14 (.A ( DP_OP_1003J1_66_5789_n55 ) 
    , .B ( DP_OP_1003J1_66_5789_n52 ) , .CI ( DP_OP_1003J1_66_5789_n14 ) 
    , .CO ( DP_OP_1003J1_66_5789_n13 ) , .S ( bajo_reg_entrada[5] ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U15 (.A ( DP_OP_1003J1_66_5789_n59 ) 
    , .B ( DP_OP_1003J1_66_5789_n56 ) , .CI ( DP_OP_1003J1_66_5789_n15 ) 
    , .CO ( DP_OP_1003J1_66_5789_n14 ) , .S ( bajo_reg_entrada[4] ) ) ;
FADDX1 DP_OP_1003J1_66_5789_U16 (.A ( DP_OP_1003J1_66_5789_n63 ) 
    , .B ( DP_OP_1003J1_66_5789_n60 ) , .CI ( DP_OP_1003J1_66_5789_n16 ) 
    , .CO ( DP_OP_1003J1_66_5789_n15 ) , .S ( bajo_reg_entrada[3] ) ) ;
FADDX1 DP_OP_1001J1_64_4995_U7 (.A ( coeficiente_b11_H_v_out[14] ) 
    , .B ( partial_2_H[14] ) , .CI ( DP_OP_1001J1_64_4995_n7 ) 
    , .CO ( DP_OP_1001J1_64_4995_n6 ) , .S ( partial_3_H[14] ) ) ;
OA221X1 U102 (.IN2 ( reloj_secuencia[4] ) , .IN4 ( reloj_secuencia[5] ) 
    , .Q ( secuencia_reloj_prioridad_salida_pre_1_ ) , .IN5 ( n1032 ) 
    , .IN1 ( n1120 ) , .IN3 ( n1120 ) ) ;
DFFASX1 sos2_reg_pila_registro_reg_7_registro_tmp_reg_0_ (.SETB ( n1659 ) 
    , .QN ( \sos2_reg/bank_registro_registros[7][0] ) 
    , .CLK ( reloj_secuencia[7] ) , .D ( n1563 ) ) ;
DFFASX1 sos2_reg_pila_registro_reg_6_registro_tmp_reg_0_ (.SETB ( n1658 ) 
    , .QN ( \sos2_reg/bank_registro_registros[6][0] ) 
    , .CLK ( reloj_secuencia[6] ) , .D ( n1563 ) ) ;
DFFASX1 sos2_reg_pila_registro_reg_5_registro_tmp_reg_0_ (.SETB ( n1658 ) 
    , .QN ( \sos2_reg/bank_registro_registros[5][0] ) 
    , .CLK ( reloj_secuencia[5] ) , .D ( n1563 ) ) ;
DFFASX1 sos2_reg_pila_registro_reg_4_registro_tmp_reg_0_ (.SETB ( n1659 ) 
    , .QN ( \sos2_reg/bank_registro_registros[4][0] ) 
    , .CLK ( reloj_secuencia[4] ) , .D ( n1563 ) ) ;
DFFASX1 sos2_reg_pila_registro_reg_3_registro_tmp_reg_0_ (.SETB ( n1650 ) 
    , .QN ( \sos2_reg/bank_registro_registros[3][0] ) 
    , .CLK ( reloj_secuencia[3] ) , .D ( n1563 ) ) ;
DFFASX1 sos2_reg_pila_registro_reg_2_registro_tmp_reg_0_ (.SETB ( n1653 ) 
    , .QN ( \sos2_reg/bank_registro_registros[2][0] ) 
    , .CLK ( reloj_secuencia[2] ) , .D ( n1563 ) ) ;
DFFASX1 sos2_reg_pila_registro_reg_1_registro_tmp_reg_0_ (.SETB ( n1652 ) 
    , .QN ( \sos2_reg/bank_registro_registros[1][0] ) 
    , .CLK ( reloj_secuencia[1] ) , .D ( n1563 ) ) ;
FADDX1 U511 (.A ( sos2_reg_entrada[12] ) , .B ( DP_OP_1002J1_65_247_n66 ) 
    , .CI ( DP_OP_1002J1_65_247_n61 ) , .CO ( DP_OP_1002J1_65_247_n58 ) 
    , .S ( DP_OP_1002J1_65_247_n59 ) ) ;
FADDX1 U510 (.A ( sos2_reg_entrada[13] ) , .B ( DP_OP_1002J1_65_247_n60 ) 
    , .CI ( DP_OP_1002J1_65_247_n55 ) , .CO ( DP_OP_1002J1_65_247_n52 ) 
    , .S ( DP_OP_1002J1_65_247_n53 ) ) ;
FADDX1 U509 (.A ( n1588 ) , .B ( DP_OP_1002J1_65_247_n54 ) 
    , .CI ( DP_OP_1002J1_65_247_n49 ) , .CO ( DP_OP_1002J1_65_247_n46 ) 
    , .S ( DP_OP_1002J1_65_247_n47 ) ) ;
INVX0 U508 (.ZN ( n1594 ) , .INP ( sos2_reg_entrada[6] ) ) ;
INVX0 U507 (.ZN ( n1595 ) , .INP ( sos2_reg_entrada[7] ) ) ;
FADDX1 U506 (.A ( sos2_reg_entrada[18] ) , .B ( sos2_reg_entrada[16] ) 
    , .CI ( sos2_reg_entrada[11] ) , .CO ( DP_OP_1002J1_65_247_n54 ) 
    , .S ( DP_OP_1002J1_65_247_n55 ) ) ;
FADDX1 U505 (.A ( sos2_reg_entrada[14] ) , .B ( sos2_reg_entrada[17] ) 
    , .CI ( sos2_reg_entrada[12] ) , .CO ( DP_OP_1002J1_65_247_n48 ) 
    , .S ( DP_OP_1002J1_65_247_n49 ) ) ;
FADDX1 U504 (.A ( sos2_reg_entrada[15] ) , .B ( sos2_reg_entrada[13] ) 
    , .CI ( n1588 ) , .CO ( DP_OP_1002J1_65_247_n42 ) 
    , .S ( DP_OP_1002J1_65_247_n43 ) ) ;
FADDX1 U519 (.A ( sos2_reg_entrada[7] ) , .B ( n1597 ) , .CI ( n1582 ) 
    , .CO ( DP_OP_1002J1_65_247_n200 ) , .S ( DP_OP_1002J1_65_247_n201 ) ) ;
FADDX1 U518 (.A ( sos2_reg_entrada[6] ) , .B ( n1596 ) , .CI ( n1581 ) 
    , .CO ( DP_OP_1002J1_65_247_n202 ) , .S ( DP_OP_1002J1_65_247_n203 ) ) ;
FADDX1 U517 (.A ( sos2_reg_entrada[11] ) , .B ( DP_OP_1002J1_65_247_n72 ) 
    , .CI ( DP_OP_1002J1_65_247_n67 ) , .CO ( DP_OP_1002J1_65_247_n64 ) 
    , .S ( DP_OP_1002J1_65_247_n65 ) ) ;
INVX0 U516 (.ZN ( n1575 ) , .INP ( DP_OP_1002J1_65_247_n261 ) ) ;
INVX0 U515 (.ZN ( n1593 ) , .INP ( sos2_reg_entrada[5] ) ) ;
FADDX1 U514 (.A ( sos2_reg_entrada[3] ) , .B ( n1593 ) , .CI ( n1595 ) 
    , .CO ( DP_OP_1002J1_65_247_n208 ) , .S ( DP_OP_1002J1_65_247_n209 ) ) ;
FADDX1 U513 (.A ( sos2_reg_entrada[4] ) , .B ( n1594 ) , .CI ( n1596 ) 
    , .CO ( DP_OP_1002J1_65_247_n206 ) , .S ( DP_OP_1002J1_65_247_n207 ) ) ;
FADDX1 U512 (.A ( sos2_reg_entrada[5] ) , .B ( n1595 ) , .CI ( n1597 ) 
    , .CO ( DP_OP_1002J1_65_247_n204 ) , .S ( DP_OP_1002J1_65_247_n205 ) ) ;
INVX0 U527 (.ZN ( n1574 ) , .INP ( DP_OP_1002J1_65_247_n262 ) ) ;
FADDX1 U526 (.A ( DP_OP_1002J1_65_247_n263 ) , .B ( DP_OP_1002J1_65_247_n35 ) 
    , .CI ( DP_OP_1002J1_65_247_n13 ) , .CO ( DP_OP_1002J1_65_247_n12 ) 
    , .S ( coeficiente_b12_H_v_out[7] ) ) ;
INVX0 U525 (.ZN ( n1573 ) , .INP ( DP_OP_1002J1_65_247_n263 ) ) ;
INVX0 U524 (.ZN ( n1572 ) , .INP ( DP_OP_1002J1_65_247_n264 ) ) ;
FADDX1 U523 (.A ( sos2_reg_entrada[16] ) , .B ( n1588 ) 
    , .CI ( DP_OP_1002J1_65_247_n32 ) , .CO ( DP_OP_1002J1_65_247_n28 ) 
    , .S ( DP_OP_1002J1_65_247_n29 ) ) ;
INVX0 U522 (.ZN ( n1592 ) , .INP ( sos2_reg_entrada[4] ) ) ;
FADDX1 U521 (.A ( sos2_reg_entrada[1] ) , .B ( n1591 ) , .CI ( n1593 ) 
    , .CO ( DP_OP_1002J1_65_247_n212 ) , .S ( DP_OP_1002J1_65_247_n213 ) ) ;
FADDX1 U520 (.A ( sos2_reg_entrada[15] ) , .B ( n1583 ) 
    , .CI ( DP_OP_1002J1_65_247_n143 ) , .CO ( DP_OP_1002J1_65_247_n141 ) 
    , .S ( DP_OP_1002J1_65_247_n142 ) ) ;
FADDX1 U535 (.A ( sos2_reg_entrada[11] ) , .B ( n1584 ) , .CI ( n1586 ) 
    , .CO ( DP_OP_1002J1_65_247_n192 ) , .S ( DP_OP_1002J1_65_247_n193 ) ) ;
FADDX1 U534 (.A ( sos2_reg_entrada[12] ) , .B ( n1585 ) , .CI ( n1560 ) 
    , .CO ( DP_OP_1002J1_65_247_n190 ) , .S ( DP_OP_1002J1_65_247_n191 ) ) ;
FADDX1 U533 (.A ( sos2_reg_entrada[13] ) , .B ( n1586 ) , .CI ( n1587 ) 
    , .CO ( DP_OP_1002J1_65_247_n188 ) , .S ( DP_OP_1002J1_65_247_n189 ) ) ;
FADDX1 U532 (.A ( sos2_reg_entrada[18] ) , .B ( n1586 ) 
    , .CI ( DP_OP_1002J1_65_247_n137 ) , .CO ( DP_OP_1002J1_65_247_n135 ) 
    , .S ( DP_OP_1002J1_65_247_n136 ) ) ;
INVX0 U531 (.ZN ( n1589 ) , .INP ( DP_OP_1002J1_65_247_n256 ) ) ;
INVX0 U530 (.ZN ( n1577 ) , .INP ( DP_OP_1002J1_65_247_n259 ) ) ;
INVX0 U529 (.ZN ( n1576 ) , .INP ( DP_OP_1002J1_65_247_n260 ) ) ;
FADDX1 U528 (.A ( DP_OP_1002J1_65_247_n261 ) , .B ( DP_OP_1002J1_65_247_n45 ) 
    , .CI ( DP_OP_1002J1_65_247_n15 ) , .CO ( DP_OP_1002J1_65_247_n14 ) 
    , .S ( coeficiente_b12_H_v_out[5] ) ) ;
AO22X1 U543 (.IN1 ( n2030 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][15] ) , .Q ( n1688 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][15] ) ) ;
AO22X1 U542 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][15] ) , .Q ( n1691 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][15] ) ) ;
INVX0 U541 (.ZN ( n1591 ) , .INP ( sos2_reg_entrada[3] ) ) ;
XOR2X1 U540 (.IN2 ( sos2_reg_entrada[0] ) , .Q ( DP_OP_1002J1_65_247_n215 ) 
    , .IN1 ( sos2_reg_entrada[2] ) ) ;
NAND2X1 U539 (.IN2 ( n1563 ) , .IN1 ( sos2_reg_entrada[2] ) 
    , .QN ( DP_OP_1002J1_65_247_n214 ) ) ;
FADDX1 U538 (.A ( sos2_reg_entrada[9] ) , .B ( n1582 ) , .CI ( n1584 ) 
    , .CO ( DP_OP_1002J1_65_247_n196 ) , .S ( DP_OP_1002J1_65_247_n197 ) ) ;
FADDX1 U537 (.A ( sos2_reg_entrada[8] ) , .B ( n1581 ) , .CI ( n1583 ) 
    , .CO ( DP_OP_1002J1_65_247_n198 ) , .S ( DP_OP_1002J1_65_247_n199 ) ) ;
FADDX1 U536 (.A ( sos2_reg_entrada[10] ) , .B ( n1583 ) , .CI ( n1585 ) 
    , .CO ( DP_OP_1002J1_65_247_n194 ) , .S ( DP_OP_1002J1_65_247_n195 ) ) ;
FADDX1 U551 (.A ( n1588 ) , .B ( n1570 ) , .CI ( DP_OP_1002J1_65_247_n24 ) 
    , .CO ( DP_OP_1002J1_65_247_n22 ) , .S ( DP_OP_1002J1_65_247_n23 ) ) ;
FADDX1 U550 (.A ( sos2_reg_entrada[14] ) , .B ( sos2_reg_entrada[16] ) 
    , .CI ( sos2_reg_entrada[18] ) , .CO ( DP_OP_1002J1_65_247_n186 ) 
    , .S ( DP_OP_1002J1_65_247_n187 ) ) ;
INVX2 U549 (.INP ( sos2_reg_entrada[15] ) , .ZN ( n1586 ) ) ;
INVX0 U548 (.ZN ( n1525 ) , .INP ( coeficiente_a11_H_in[12] ) ) ;
AO22X1 U547 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][7] ) , .Q ( n1728 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][7] ) ) ;
AO22X1 U546 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][7] ) , .Q ( n1731 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][7] ) ) ;
AO22X1 U545 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][8] ) , .Q ( n1732 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][8] ) ) ;
AO22X1 U544 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][8] ) , .Q ( n1735 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][8] ) ) ;
FADDX1 U559 (.A ( coeficiente_a11_H_in[15] ) , .B ( coeficiente_a11_H_in[17] ) 
    , .CI ( coeficiente_b12_H_v_out[6] ) , .CO ( DP_OP_1001J1_64_4995_n96 ) 
    , .S ( DP_OP_1001J1_64_4995_n97 ) ) ;
FADDX1 U558 (.A ( coeficiente_b12_H_v_out[7] ) , .B ( n1528 ) , .CI ( n1529 ) 
    , .CO ( DP_OP_1001J1_64_4995_n90 ) , .S ( DP_OP_1001J1_64_4995_n91 ) ) ;
FADDX1 U557 (.A ( DP_OP_1002J1_65_247_n264 ) , .B ( DP_OP_1002J1_65_247_n31 ) 
    , .CI ( DP_OP_1002J1_65_247_n12 ) , .CO ( DP_OP_1002J1_65_247_n11 ) 
    , .S ( coeficiente_b12_H_v_out[8] ) ) ;
AO22X1 U556 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][17] ) , .Q ( n1696 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][17] ) ) ;
AO22X1 U555 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][17] ) , .Q ( n1699 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][17] ) ) ;
INVX0 U554 (.ZN ( n1571 ) , .INP ( DP_OP_1002J1_65_247_n265 ) ) ;
FADDX1 U553 (.A ( sos2_reg_entrada[17] ) , .B ( DP_OP_1002J1_65_247_n28 ) 
    , .CI ( DP_OP_1002J1_65_247_n26 ) , .CO ( DP_OP_1002J1_65_247_n24 ) 
    , .S ( DP_OP_1002J1_65_247_n25 ) ) ;
INVX0 U552 (.ZN ( n1570 ) , .INP ( DP_OP_1002J1_65_247_n266 ) ) ;
AO22X1 U567 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][12] ) , .Q ( n1679 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][12] ) ) ;
INVX0 U566 (.ZN ( n1579 ) , .INP ( DP_OP_1002J1_65_247_n257 ) ) ;
INVX0 U565 (.ZN ( n1523 ) , .INP ( coeficiente_a11_H_in[10] ) ) ;
INVX0 U564 (.ZN ( n1524 ) , .INP ( coeficiente_a11_H_in[11] ) ) ;
INVX0 U563 (.ZN ( n1578 ) , .INP ( DP_OP_1002J1_65_247_n258 ) ) ;
AO22X1 U562 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][18] ) , .Q ( n1700 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][18] ) ) ;
AO22X1 U561 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][18] ) , .Q ( n1703 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][18] ) ) ;
FADDX1 U560 (.A ( coeficiente_a11_H_in[14] ) , .B ( coeficiente_a11_H_in[16] ) 
    , .CI ( coeficiente_b12_H_v_out[5] ) , .CO ( DP_OP_1001J1_64_4995_n102 ) 
    , .S ( DP_OP_1001J1_64_4995_n103 ) ) ;
INVX2 U575 (.INP ( sos2_reg_entrada[16] ) , .ZN ( n1560 ) ) ;
FADDX1 U574 (.A ( sos2_reg_entrada[16] ) , .B ( n1588 ) 
    , .CI ( DP_OP_1002J1_65_247_n135 ) , .CO ( DP_OP_1002J1_65_247_n133 ) 
    , .S ( DP_OP_1002J1_65_247_n134 ) ) ;
FADDX1 U573 (.A ( sos2_reg_entrada[7] ) , .B ( sos2_reg_entrada[12] ) 
    , .CI ( sos2_reg_entrada[9] ) , .CO ( DP_OP_1002J1_65_247_n74 ) 
    , .S ( DP_OP_1002J1_65_247_n75 ) ) ;
AO22X1 U572 (.IN1 ( n2030 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][14] ) , .Q ( n1684 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][14] ) ) ;
AO22X1 U571 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][14] ) , .Q ( n1687 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][14] ) ) ;
AO22X1 U570 (.IN1 ( n2030 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][10] ) , .Q ( n1668 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][10] ) ) ;
AO22X1 U569 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][10] ) , .Q ( n1671 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][10] ) ) ;
AO22X1 U568 (.IN1 ( n2030 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][12] ) , .Q ( n1676 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][12] ) ) ;
INVX0 U583 (.ZN ( n1555 ) , .INP ( coeficiente_b11_L_v_out[15] ) ) ;
INVX0 U582 (.ZN ( n1556 ) , .INP ( coeficiente_b11_L_v_out[16] ) ) ;
INVX0 U581 (.ZN ( n1552 ) , .INP ( coeficiente_b11_L_v_out[12] ) ) ;
FADDX1 U580 (.A ( coeficiente_b12_L_v_out[3] ) 
    , .B ( coeficiente_b11_L_v_out[14] ) , .CI ( n1552 ) 
    , .CO ( DP_OP_1001J1_64_4995_n261 ) , .S ( DP_OP_1001J1_64_4995_n262 ) ) ;
INVX0 U579 (.ZN ( n1557 ) , .INP ( coeficiente_b11_L_v_out[17] ) ) ;
FADDX1 U578 (.A ( coeficiente_b12_L_v_out[4] ) 
    , .B ( coeficiente_b11_L_v_out[15] ) , .CI ( n1553 ) 
    , .CO ( DP_OP_1001J1_64_4995_n255 ) , .S ( DP_OP_1001J1_64_4995_n256 ) ) ;
FADDX1 U577 (.A ( coeficiente_b11_L_v_out[14] ) 
    , .B ( coeficiente_b11_L_v_out[16] ) , .CI ( coeficiente_b12_L_v_out[5] ) 
    , .CO ( DP_OP_1001J1_64_4995_n249 ) , .S ( DP_OP_1001J1_64_4995_n250 ) ) ;
FADDX1 U576 (.A ( coeficiente_b11_L_v_out[15] ) 
    , .B ( coeficiente_b11_L_v_out[17] ) , .CI ( coeficiente_b12_L_v_out[6] ) 
    , .CO ( DP_OP_1001J1_64_4995_n243 ) , .S ( DP_OP_1001J1_64_4995_n244 ) ) ;
INVX0 U591 (.ZN ( n1530 ) , .INP ( coeficiente_a11_H_in[17] ) ) ;
INVX0 U590 (.ZN ( n1531 ) , .INP ( coeficiente_a11_H_in[18] ) ) ;
INVX0 U589 (.ZN ( n1528 ) , .INP ( coeficiente_a11_H_in[15] ) ) ;
AO22X1 U588 (.IN1 ( n1643 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][16] ) , .Q ( n1692 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][16] ) ) ;
AO22X1 U587 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][16] ) , .Q ( n1695 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][16] ) ) ;
INVX0 U586 (.ZN ( n1590 ) , .INP ( sos2_reg_entrada[1] ) ) ;
AO22X1 U585 (.IN1 ( n1643 ) , .IN3 ( n1640 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][12] ) , .Q ( n1828 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][12] ) ) ;
AO22X1 U584 (.IN1 ( n2028 ) , .IN3 ( n1634 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][12] ) , .Q ( n1829 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][12] ) ) ;
AO22X1 U599 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][4] ) , .Q ( n1716 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][4] ) ) ;
AO22X1 U598 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][4] ) , .Q ( n1719 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][4] ) ) ;
AO22X1 U597 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][6] ) , .Q ( n1724 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][6] ) ) ;
AO22X1 U596 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][6] ) , .Q ( n1727 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][6] ) ) ;
AO22X1 U595 (.IN1 ( n2030 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][3] ) , .Q ( n1712 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][3] ) ) ;
AO22X1 U594 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][3] ) , .Q ( n1715 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][3] ) ) ;
INVX0 U593 (.ZN ( n1615 ) , .INP ( partial_3_H[15] ) ) ;
INVX0 U592 (.ZN ( n1620 ) , .INP ( partial_3_H[10] ) ) ;
AO22X1 U607 (.IN1 ( n1643 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][15] ) , .Q ( n1840 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][15] ) ) ;
AO22X1 U606 (.IN1 ( n2030 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][2] ) , .Q ( n1708 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][2] ) ) ;
AO22X1 U605 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][2] ) , .Q ( n1711 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][2] ) ) ;
AO22X1 U604 (.IN1 ( n2030 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][1] ) , .Q ( n1704 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][1] ) ) ;
AO22X1 U603 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][1] ) , .Q ( n1707 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][1] ) ) ;
INVX0 U602 (.ZN ( n1506 ) , .INP ( coeficiente_b11_H_v_out[0] ) ) ;
AO22X1 U601 (.IN1 ( n1641 ) , .IN3 ( n1639 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][0] ) , .Q ( n1664 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][0] ) ) ;
AO22X1 U600 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][0] ) , .Q ( n1667 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][0] ) ) ;
AO22X1 U615 (.IN1 ( n1641 ) , .IN3 ( n1640 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][8] ) , .Q ( n1884 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][8] ) ) ;
AO22X1 U614 (.IN1 ( n2028 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][8] ) , .Q ( n1885 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][8] ) ) ;
INVX0 U613 (.ZN ( n1604 ) , .INP ( partial_3_L[13] ) ) ;
INVX0 U612 (.ZN ( n1603 ) , .INP ( partial_3_L[14] ) ) ;
AO22X1 U611 (.IN1 ( n1643 ) , .IN3 ( n1640 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][18] ) , .Q ( n1852 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][18] ) ) ;
AO22X1 U610 (.IN1 ( n1637 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][18] ) , .Q ( n1853 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][18] ) ) ;
AO22X1 U609 (.IN1 ( n1643 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][14] ) , .Q ( n1836 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][14] ) ) ;
AO22X1 U608 (.IN1 ( n1637 ) , .IN3 ( n1634 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][14] ) , .Q ( n1837 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][14] ) ) ;
AO22X1 U623 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( bank_registro_registros[78] ) , .Q ( n1963 ) 
    , .IN4 ( bank_registro_registros[96] ) ) ;
AO22X1 U622 (.IN1 ( n2030 ) , .IN3 ( n2029 ) 
    , .IN2 ( bank_registro_registros[61] ) , .Q ( n1964 ) 
    , .IN4 ( bank_registro_registros[43] ) ) ;
AO22X1 U621 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( bank_registro_registros[79] ) , .Q ( n1967 ) 
    , .IN4 ( bank_registro_registros[97] ) ) ;
AO22X1 U620 (.IN1 ( n2030 ) , .IN3 ( n1640 ) 
    , .IN2 ( bank_registro_registros[62] ) , .Q ( n1896 ) 
    , .IN4 ( bank_registro_registros[44] ) ) ;
AO22X1 U619 (.IN1 ( n2028 ) , .IN3 ( n1634 ) 
    , .IN2 ( bank_registro_registros[10] ) , .Q ( n1897 ) 
    , .IN4 ( bank_registro_registros[26] ) ) ;
INVX0 U618 (.ZN ( n1536 ) , .INP ( coeficiente_a22_in[14] ) ) ;
AO22X1 U617 (.IN1 ( n1642 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][10] ) , .Q ( n1820 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][10] ) ) ;
AO22X1 U616 (.IN1 ( n2028 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][10] ) , .Q ( n1821 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][10] ) ) ;
AO22X1 U631 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( bank_registro_registros[76] ) , .Q ( n1955 ) 
    , .IN4 ( bank_registro_registros[94] ) ) ;
FADDX1 U630 (.A ( coeficiente_a22_in[10] ) , .B ( n1539 ) , .CI ( n1587 ) 
    , .CO ( DP_OP_1001J1_64_4995_n408 ) , .S ( DP_OP_1001J1_64_4995_n409 ) ) ;
AO22X1 U629 (.IN1 ( n1642 ) , .IN3 ( n2029 ) 
    , .IN2 ( bank_registro_registros[59] ) , .Q ( n1956 ) 
    , .IN4 ( bank_registro_registros[41] ) ) ;
AO22X1 U628 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( bank_registro_registros[77] ) , .Q ( n1959 ) 
    , .IN4 ( bank_registro_registros[95] ) ) ;
INVX0 U627 (.ZN ( n1548 ) , .INP ( coeficiente_a22_in[8] ) ) ;
INVX0 U626 (.ZN ( n1549 ) , .INP ( coeficiente_a22_in[9] ) ) ;
FADDX1 U625 (.A ( n1586 ) , .B ( n1549 ) , .CI ( n1560 ) 
    , .CO ( DP_OP_1001J1_64_4995_n384 ) , .S ( DP_OP_1001J1_64_4995_n385 ) ) ;
AO22X1 U624 (.IN1 ( n1642 ) , .IN3 ( n2029 ) 
    , .IN2 ( bank_registro_registros[60] ) , .Q ( n1960 ) 
    , .IN4 ( bank_registro_registros[42] ) ) ;
AO22X1 U639 (.IN1 ( n1642 ) , .IN3 ( n1640 ) 
    , .IN2 ( bank_registro_registros[56] ) , .Q ( n1944 ) 
    , .IN4 ( bank_registro_registros[38] ) ) ;
AO22X1 U638 (.IN1 ( n1637 ) , .IN3 ( n2027 ) 
    , .IN2 ( bank_registro_registros[4] ) , .Q ( n1945 ) 
    , .IN4 ( bank_registro_registros[20] ) ) ;
FADDX1 U637 (.A ( n1538 ) , .B ( n1540 ) , .CI ( sos2_reg_entrada[18] ) 
    , .CO ( DP_OP_1001J1_64_4995_n420 ) , .S ( DP_OP_1001J1_64_4995_n421 ) ) ;
AO22X1 U636 (.IN1 ( n1642 ) , .IN3 ( n2029 ) 
    , .IN2 ( bank_registro_registros[57] ) , .Q ( n1948 ) 
    , .IN4 ( bank_registro_registros[39] ) ) ;
AO22X1 U635 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( bank_registro_registros[75] ) , .Q ( n1951 ) 
    , .IN4 ( bank_registro_registros[93] ) ) ;
INVX0 U634 (.ZN ( n1546 ) , .INP ( coeficiente_a22_in[6] ) ) ;
INVX0 U633 (.ZN ( n1547 ) , .INP ( coeficiente_a22_in[7] ) ) ;
AO22X1 U632 (.IN1 ( n1642 ) , .IN3 ( n2029 ) 
    , .IN2 ( bank_registro_registros[58] ) , .Q ( n1952 ) 
    , .IN4 ( bank_registro_registros[40] ) ) ;
INVX0 U647 (.ZN ( n1537 ) , .INP ( coeficiente_a22_in[15] ) ) ;
AO22X1 U646 (.IN1 ( n1642 ) , .IN3 ( n2029 ) 
    , .IN2 ( bank_registro_registros[54] ) , .Q ( n1936 ) 
    , .IN4 ( bank_registro_registros[36] ) ) ;
AO22X1 U645 (.IN1 ( n2028 ) , .IN3 ( n2027 ) 
    , .IN2 ( bank_registro_registros[2] ) , .Q ( n1937 ) 
    , .IN4 ( bank_registro_registros[18] ) ) ;
INVX0 U644 (.ZN ( n1581 ) , .INP ( sos2_reg_entrada[10] ) ) ;
INVX0 U643 (.ZN ( n1544 ) , .INP ( coeficiente_a22_in[4] ) ) ;
AO22X1 U642 (.IN1 ( n1642 ) , .IN3 ( n2029 ) 
    , .IN2 ( bank_registro_registros[55] ) , .Q ( n1940 ) 
    , .IN4 ( bank_registro_registros[37] ) ) ;
AO22X1 U641 (.IN1 ( n1637 ) , .IN3 ( n1634 ) 
    , .IN2 ( bank_registro_registros[3] ) , .Q ( n1941 ) 
    , .IN4 ( bank_registro_registros[19] ) ) ;
INVX0 U640 (.ZN ( n1545 ) , .INP ( coeficiente_a22_in[5] ) ) ;
FADDX1 U655 (.A ( sos2_reg_entrada[15] ) , .B ( sos2_reg_entrada[17] ) 
    , .CI ( n1560 ) , .CO ( DP_OP_1002J1_65_247_n184 ) 
    , .S ( DP_OP_1002J1_65_247_n185 ) ) ;
INVX0 U654 (.ZN ( n1534 ) , .INP ( coeficiente_a22_in[12] ) ) ;
INVX0 U653 (.ZN ( n1597 ) , .INP ( sos2_reg_entrada[9] ) ) ;
INVX0 U652 (.ZN ( n1583 ) , .INP ( sos2_reg_entrada[12] ) ) ;
INVX2 U651 (.INP ( sos2_reg_entrada[13] ) , .ZN ( n1584 ) ) ;
INVX2 U650 (.INP ( sos2_reg_entrada[14] ) , .ZN ( n1585 ) ) ;
INVX0 U649 (.ZN ( n1535 ) , .INP ( coeficiente_a22_in[13] ) ) ;
FADDX1 U648 (.A ( coeficiente_a22_in[6] ) , .B ( coeficiente_a22_in[8] ) 
    , .CI ( n1586 ) , .CO ( DP_OP_1001J1_64_4995_n464 ) 
    , .S ( DP_OP_1001J1_64_4995_n465 ) ) ;
FADDX1 U663 (.A ( n1531 ) , .B ( DP_OP_1001J1_64_4995_n96 ) 
    , .CI ( DP_OP_1001J1_64_4995_n91 ) , .CO ( DP_OP_1001J1_64_4995_n88 ) 
    , .S ( DP_OP_1001J1_64_4995_n89 ) ) ;
FADDX1 U662 (.A ( coeficiente_b12_H_v_out[9] ) , .B ( n1530 ) 
    , .CI ( coeficiente_a11_H_in[18] ) , .CO ( DP_OP_1001J1_64_4995_n80 ) 
    , .S ( DP_OP_1001J1_64_4995_n81 ) ) ;
FADDX1 U661 (.A ( DP_OP_1002J1_65_247_n266 ) , .B ( DP_OP_1002J1_65_247_n25 ) 
    , .CI ( DP_OP_1002J1_65_247_n10 ) , .CO ( DP_OP_1002J1_65_247_n9 ) 
    , .S ( coeficiente_b12_H_v_out[10] ) ) ;
INVX0 U660 (.ZN ( n1569 ) , .INP ( DP_OP_1002J1_65_247_n267 ) ) ;
INVX0 U659 (.ZN ( n1568 ) , .INP ( DP_OP_1002J1_65_247_n268 ) ) ;
INVX0 U658 (.ZN ( n1567 ) , .INP ( DP_OP_1002J1_65_247_n269 ) ) ;
INVX0 U657 (.ZN ( n1566 ) , .INP ( DP_OP_1002J1_65_247_n270 ) ) ;
INVX0 U656 (.ZN ( n1565 ) , .INP ( DP_OP_1002J1_65_247_n271 ) ) ;
AO22X1 U671 (.IN1 ( n2030 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][11] ) , .Q ( n1672 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][11] ) ) ;
AO22X1 U670 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][11] ) , .Q ( n1675 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][11] ) ) ;
INVX0 U669 (.ZN ( n1527 ) , .INP ( coeficiente_a11_H_in[14] ) ) ;
FADDX1 U668 (.A ( n1528 ) , .B ( n1523 ) , .CI ( DP_OP_1001J1_64_4995_n124 ) 
    , .CO ( DP_OP_1001J1_64_4995_n118 ) , .S ( DP_OP_1001J1_64_4995_n119 ) ) ;
FADDX1 U667 (.A ( n1529 ) , .B ( DP_OP_1001J1_64_4995_n120 ) 
    , .CI ( DP_OP_1001J1_64_4995_n115 ) , .CO ( DP_OP_1001J1_64_4995_n112 ) 
    , .S ( DP_OP_1001J1_64_4995_n113 ) ) ;
FADDX1 U666 (.A ( n1530 ) , .B ( DP_OP_1001J1_64_4995_n114 ) 
    , .CI ( DP_OP_1001J1_64_4995_n109 ) , .CO ( DP_OP_1001J1_64_4995_n106 ) 
    , .S ( DP_OP_1001J1_64_4995_n107 ) ) ;
FADDX1 U665 (.A ( coeficiente_a11_H_in[18] ) 
    , .B ( DP_OP_1001J1_64_4995_n108 ) , .CI ( DP_OP_1001J1_64_4995_n103 ) 
    , .CO ( DP_OP_1001J1_64_4995_n100 ) , .S ( DP_OP_1001J1_64_4995_n101 ) ) ;
FADDX1 U664 (.A ( n1527 ) , .B ( DP_OP_1001J1_64_4995_n102 ) 
    , .CI ( DP_OP_1001J1_64_4995_n97 ) , .CO ( DP_OP_1001J1_64_4995_n94 ) 
    , .S ( DP_OP_1001J1_64_4995_n95 ) ) ;
FADDX1 U679 (.A ( n1580 ) , .B ( DP_OP_1002J1_65_247_n272 ) 
    , .CI ( DP_OP_1002J1_65_247_n101 ) , .CO ( DP_OP_1002J1_65_247_n100 ) 
    , .S ( coeficiente_b12_L_v_out[16] ) ) ;
FADDX1 U678 (.A ( sos2_reg_entrada[16] ) , .B ( n1587 ) 
    , .CI ( sos2_reg_entrada[18] ) , .CO ( DP_OP_1002J1_65_247_n182 ) 
    , .S ( DP_OP_1002J1_65_247_n183 ) ) ;
INVX2 U677 (.INP ( DP_OP_1002J1_65_247_n127 ) , .ZN ( n1580 ) ) ;
FADDX1 U676 (.A ( sos2_reg_entrada[17] ) , .B ( n1560 ) 
    , .CI ( DP_OP_1002J1_65_247_n133 ) , .CO ( DP_OP_1002J1_65_247_n131 ) 
    , .S ( DP_OP_1002J1_65_247_n132 ) ) ;
AO22X1 U675 (.IN1 ( n2030 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][13] ) , .Q ( n1680 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][13] ) ) ;
AO22X1 U674 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][13] ) , .Q ( n1683 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][13] ) ) ;
AO22X1 U673 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][9] ) , .Q ( n1736 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][9] ) ) ;
AO22X1 U672 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][9] ) , .Q ( n1739 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][9] ) ) ;
FADDX1 U687 (.A ( n1580 ) , .B ( DP_OP_1002J1_65_247_n268 ) 
    , .CI ( DP_OP_1002J1_65_247_n105 ) , .CO ( DP_OP_1002J1_65_247_n104 ) 
    , .S ( coeficiente_b12_L_v_out[12] ) ) ;
FADDX1 U686 (.A ( n1580 ) , .B ( DP_OP_1002J1_65_247_n269 ) 
    , .CI ( DP_OP_1002J1_65_247_n104 ) , .CO ( DP_OP_1002J1_65_247_n103 ) 
    , .S ( coeficiente_b12_L_v_out[13] ) ) ;
AO22X1 U685 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][14] ) , .Q ( n1760 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][14] ) ) ;
AO22X1 U684 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][14] ) , .Q ( n1763 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][14] ) ) ;
FADDX1 U683 (.A ( n1580 ) , .B ( DP_OP_1002J1_65_247_n270 ) 
    , .CI ( DP_OP_1002J1_65_247_n103 ) , .CO ( DP_OP_1002J1_65_247_n102 ) 
    , .S ( coeficiente_b12_L_v_out[14] ) ) ;
AO22X1 U682 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][15] ) , .Q ( n1764 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][15] ) ) ;
AO22X1 U681 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][15] ) , .Q ( n1767 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][15] ) ) ;
FADDX1 U680 (.A ( n1580 ) , .B ( DP_OP_1002J1_65_247_n271 ) 
    , .CI ( DP_OP_1002J1_65_247_n102 ) , .CO ( DP_OP_1002J1_65_247_n101 ) 
    , .S ( coeficiente_b12_L_v_out[15] ) ) ;
AO22X1 U695 (.IN1 ( n1641 ) , .IN3 ( n1640 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][9] ) , .Q ( n1812 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][9] ) ) ;
AO22X1 U694 (.IN1 ( n2028 ) , .IN3 ( n1634 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][9] ) , .Q ( n1813 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][9] ) ) ;
AO22X1 U693 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][10] ) , .Q ( n1744 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][10] ) ) ;
AO22X1 U692 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][10] ) , .Q ( n1747 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][10] ) ) ;
AO22X1 U691 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][11] ) , .Q ( n1748 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][11] ) ) ;
AO22X1 U690 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][11] ) , .Q ( n1751 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][11] ) ) ;
AO22X1 U689 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][12] ) , .Q ( n1752 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][12] ) ) ;
AO22X1 U688 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][12] ) , .Q ( n1755 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][12] ) ) ;
AO22X1 U703 (.IN1 ( n2028 ) , .IN3 ( n1634 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][5] ) , .Q ( n1797 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][5] ) ) ;
FADDX1 U702 (.A ( coeficiente_b11_L_v_out[18] ) 
    , .B ( DP_OP_1001J1_64_4995_n255 ) , .CI ( DP_OP_1001J1_64_4995_n250 ) 
    , .CO ( DP_OP_1001J1_64_4995_n247 ) , .S ( DP_OP_1001J1_64_4995_n248 ) ) ;
AO22X1 U701 (.IN1 ( n1642 ) , .IN3 ( n1640 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][7] ) , .Q ( n1804 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][7] ) ) ;
AO22X1 U700 (.IN1 ( n2028 ) , .IN3 ( n1633 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][7] ) , .Q ( n1805 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][7] ) ) ;
INVX0 U699 (.ZN ( n1558 ) , .INP ( coeficiente_b11_L_v_out[18] ) ) ;
AO22X1 U698 (.IN1 ( n1644 ) , .IN3 ( n1640 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][8] ) , .Q ( n1808 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][8] ) ) ;
AO22X1 U697 (.IN1 ( n2028 ) , .IN3 ( n1634 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][8] ) , .Q ( n1809 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][8] ) ) ;
FADDX1 U696 (.A ( coeficiente_b12_L_v_out[8] ) 
    , .B ( coeficiente_b11_L_v_out[17] ) , .CI ( DP_OP_1001J1_64_4995_n237 ) 
    , .CO ( DP_OP_1001J1_64_4995_n231 ) , .S ( DP_OP_1001J1_64_4995_n232 ) ) ;
INVX0 U711 (.ZN ( n1554 ) , .INP ( coeficiente_b11_L_v_out[14] ) ) ;
AO22X1 U710 (.IN1 ( n1641 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][2] ) , .Q ( n1784 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][2] ) ) ;
AO22X1 U709 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][2] ) , .Q ( n1787 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][2] ) ) ;
INVX0 U708 (.ZN ( n1550 ) , .INP ( coeficiente_b11_L_v_out[10] ) ) ;
INVX0 U707 (.ZN ( n1551 ) , .INP ( coeficiente_b11_L_v_out[11] ) ) ;
AO22X1 U706 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][3] ) , .Q ( n1788 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][3] ) ) ;
AO22X1 U705 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][3] ) , .Q ( n1791 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][3] ) ) ;
AO22X1 U704 (.IN1 ( n1643 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][5] ) , .Q ( n1796 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][5] ) ) ;
FADDX1 U719 (.A ( partial_3_H[10] ) , .B ( partial_3_H[13] ) , .CI ( n1615 ) 
    , .CO ( DP_OP_1004J1_67_3033_n41 ) , .S ( DP_OP_1004J1_67_3033_n42 ) ) ;
FADDX1 U718 (.A ( partial_3_H[11] ) , .B ( partial_3_H[14] ) , .CI ( n1614 ) 
    , .CO ( DP_OP_1004J1_67_3033_n37 ) , .S ( DP_OP_1004J1_67_3033_n38 ) ) ;
FADDX1 U717 (.A ( partial_3_H[12] ) , .B ( partial_3_H[15] ) , .CI ( n1613 ) 
    , .CO ( DP_OP_1004J1_67_3033_n33 ) , .S ( DP_OP_1004J1_67_3033_n34 ) ) ;
INVX0 U716 (.ZN ( n1529 ) , .INP ( coeficiente_a11_H_in[16] ) ) ;
AO22X1 U715 (.IN1 ( n1643 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][13] ) , .Q ( n1832 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][13] ) ) ;
AO22X1 U714 (.IN1 ( n2028 ) , .IN3 ( n1634 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][13] ) , .Q ( n1833 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][13] ) ) ;
AO22X1 U713 (.IN1 ( n1643 ) , .IN3 ( n1640 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][9] ) , .Q ( n1888 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][9] ) ) ;
AO22X1 U712 (.IN1 ( n2028 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][9] ) , .Q ( n1889 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][9] ) ) ;
INVX0 U727 (.ZN ( n1616 ) , .INP ( partial_3_H[14] ) ) ;
INVX0 U726 (.ZN ( n1622 ) , .INP ( partial_3_H[8] ) ) ;
INVX0 U725 (.ZN ( n1618 ) , .INP ( partial_3_H[12] ) ) ;
INVX0 U724 (.ZN ( n1621 ) , .INP ( partial_3_H[9] ) ) ;
FADDX1 U723 (.A ( partial_3_H[5] ) , .B ( n1620 ) , .CI ( n1616 ) 
    , .CO ( DP_OP_1004J1_67_3033_n71 ) , .S ( DP_OP_1004J1_67_3033_n72 ) ) ;
FADDX1 U722 (.A ( partial_3_H[6] ) , .B ( n1619 ) , .CI ( n1615 ) 
    , .CO ( DP_OP_1004J1_67_3033_n65 ) , .S ( DP_OP_1004J1_67_3033_n66 ) ) ;
FADDX1 U721 (.A ( n1618 ) , .B ( partial_3_H[18] ) 
    , .CI ( DP_OP_1004J1_67_3033_n65 ) , .CO ( DP_OP_1004J1_67_3033_n57 ) 
    , .S ( DP_OP_1004J1_67_3033_n58 ) ) ;
FADDX1 U720 (.A ( n1617 ) , .B ( n1614 ) , .CI ( DP_OP_1004J1_67_3033_n59 ) 
    , .CO ( DP_OP_1004J1_67_3033_n51 ) , .S ( DP_OP_1004J1_67_3033_n52 ) ) ;
AO22X1 U735 (.IN1 ( n1643 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][16] ) , .Q ( n1844 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][16] ) ) ;
AO22X1 U734 (.IN1 ( n1637 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][16] ) , .Q ( n1845 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][16] ) ) ;
AO22X1 U733 (.IN1 ( n1643 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][17] ) , .Q ( n1848 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][17] ) ) ;
AO22X1 U732 (.IN1 ( n1637 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][17] ) , .Q ( n1849 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][17] ) ) ;
INVX0 U731 (.ZN ( n1623 ) , .INP ( partial_3_H[7] ) ) ;
INVX0 U730 (.ZN ( n1619 ) , .INP ( partial_3_H[11] ) ) ;
AO22X1 U729 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[3][5] ) , .Q ( n1720 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[2][5] ) ) ;
AO22X1 U728 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[4][5] ) , .Q ( n1723 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[5][5] ) ) ;
FADDX1 U743 (.A ( partial_3_L[14] ) , .B ( partial_3_L[6] ) , .CI ( n1606 ) 
    , .CO ( DP_OP_1003J1_66_5789_n57 ) , .S ( DP_OP_1003J1_66_5789_n58 ) ) ;
INVX0 U742 (.ZN ( n1608 ) , .INP ( partial_3_L[9] ) ) ;
INVX0 U741 (.ZN ( n1607 ) , .INP ( partial_3_L[10] ) ) ;
INVX0 U740 (.ZN ( n1605 ) , .INP ( partial_3_L[12] ) ) ;
FADDX1 U739 (.A ( partial_3_L[11] ) , .B ( partial_3_L[16] ) , .CI ( n1603 ) 
    , .CO ( DP_OP_1003J1_66_5789_n37 ) , .S ( DP_OP_1003J1_66_5789_n38 ) ) ;
INVX0 U738 (.ZN ( n1602 ) , .INP ( partial_3_L[15] ) ) ;
XOR3X1 U737 (.Q ( partial_3_L[18] ) , .IN2 ( partial_2_L[18] ) 
    , .IN1 ( coeficiente_b11_L_v_out[18] ) , .IN3 ( DP_OP_1001J1_64_4995_n150 ) ) ;
FADDX1 U736 (.A ( partial_3_L[13] ) , .B ( n1600 ) , .CI ( n1601 ) 
    , .CO ( DP_OP_1003J1_66_5789_n29 ) , .S ( DP_OP_1003J1_66_5789_n30 ) ) ;
AO22X1 U751 (.IN1 ( n1637 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][7] ) , .Q ( n1881 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][7] ) ) ;
AO22X1 U750 (.IN1 ( n1643 ) , .IN3 ( n1640 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][4] ) , .Q ( n1868 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][4] ) ) ;
AO22X1 U749 (.IN1 ( n1637 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][4] ) , .Q ( n1869 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][4] ) ) ;
INVX0 U748 (.ZN ( n1609 ) , .INP ( partial_3_L[8] ) ) ;
AO22X1 U747 (.IN1 ( n1643 ) , .IN3 ( n1640 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][6] ) , .Q ( n1876 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][6] ) ) ;
AO22X1 U746 (.IN1 ( n1637 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][6] ) , .Q ( n1877 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][6] ) ) ;
AO22X1 U745 (.IN1 ( n1641 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][11] ) , .Q ( n1824 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][11] ) ) ;
AO22X1 U744 (.IN1 ( n2028 ) , .IN3 ( n1634 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][11] ) , .Q ( n1825 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][11] ) ) ;
INVX0 U759 (.ZN ( n1470 ) , .INP ( n2029 ) ) ;
AO22X1 U758 (.IN1 ( n1643 ) , .IN3 ( n2029 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][0] ) , .Q ( n1816 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][0] ) ) ;
AO22X1 U757 (.IN1 ( n1637 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][0] ) , .Q ( n1817 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][0] ) ) ;
AO22X1 U756 (.IN1 ( n1643 ) , .IN3 ( n1640 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][1] ) , .Q ( n1856 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][1] ) ) ;
AO22X1 U755 (.IN1 ( n1637 ) , .IN3 ( n1634 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][1] ) , .Q ( n1857 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][1] ) ) ;
AO22X1 U754 (.IN1 ( n1643 ) , .IN3 ( n1640 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][2] ) , .Q ( n1860 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][2] ) ) ;
AO22X1 U753 (.IN1 ( n1637 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][2] ) , .Q ( n1861 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][2] ) ) ;
AO22X1 U752 (.IN1 ( n2030 ) , .IN3 ( n1640 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][7] ) , .Q ( n1880 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][7] ) ) ;
INVX0 U767 (.ZN ( n1644 ) , .INP ( n1645 ) ) ;
AO22X1 U766 (.IN1 ( n1642 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][17] ) , .Q ( n1772 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][17] ) ) ;
AO22X1 U765 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][17] ) , .Q ( n1775 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][17] ) ) ;
INVX0 U764 (.ZN ( n1538 ) , .INP ( coeficiente_a22_in[16] ) ) ;
AO22X1 U763 (.IN1 ( n1641 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][18] ) , .Q ( n1776 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][18] ) ) ;
AO22X1 U762 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][18] ) , .Q ( n1779 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][18] ) ) ;
INVX0 U761 (.ZN ( n1539 ) , .INP ( coeficiente_a22_in[17] ) ) ;
INVX0 U760 (.ZN ( n1472 ) , .INP ( n2026 ) ) ;
AO22X1 U775 (.IN1 ( n2030 ) , .IN3 ( n2029 ) 
    , .IN2 ( bank_registro_registros[65] ) , .Q ( n1908 ) 
    , .IN4 ( bank_registro_registros[47] ) ) ;
AO22X1 U774 (.IN1 ( n2028 ) , .IN3 ( n2027 ) 
    , .IN2 ( bank_registro_registros[13] ) , .Q ( n1909 ) 
    , .IN4 ( bank_registro_registros[29] ) ) ;
FADDX1 U773 (.A ( coeficiente_a22_in[17] ) , .B ( coeficiente_a22_in[14] ) 
    , .CI ( in_reg_salida_v[13] ) , .CO ( DP_OP_1001J1_64_4995_n348 ) 
    , .S ( DP_OP_1001J1_64_4995_n349 ) ) ;
AO22X1 U772 (.IN1 ( n2030 ) , .IN3 ( n1640 ) 
    , .IN2 ( bank_registro_registros[66] ) , .Q ( n1912 ) 
    , .IN4 ( bank_registro_registros[48] ) ) ;
AO22X1 U771 (.IN1 ( n2028 ) , .IN3 ( n2027 ) 
    , .IN2 ( bank_registro_registros[14] ) , .Q ( n1913 ) 
    , .IN4 ( bank_registro_registros[30] ) ) ;
INVX0 U770 (.ZN ( n1540 ) , .INP ( coeficiente_a22_in[18] ) ) ;
AO22X1 U769 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][16] ) , .Q ( n1768 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][16] ) ) ;
AO22X1 U768 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][16] ) , .Q ( n1771 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][16] ) ) ;
INVX0 U783 (.ZN ( n1532 ) , .INP ( coeficiente_a22_in[10] ) ) ;
FADDX1 U782 (.A ( coeficiente_a22_in[13] ) , .B ( n1532 ) 
    , .CI ( DP_OP_1001J1_64_4995_n386 ) , .CO ( DP_OP_1001J1_64_4995_n374 ) 
    , .S ( DP_OP_1001J1_64_4995_n375 ) ) ;
FADDX1 U781 (.A ( coeficiente_a22_in[15] ) , .B ( DP_OP_1001J1_64_4995_n368 ) 
    , .CI ( DP_OP_1001J1_64_4995_n366 ) , .CO ( DP_OP_1001J1_64_4995_n358 ) 
    , .S ( DP_OP_1001J1_64_4995_n359 ) ) ;
AO22X1 U780 (.IN1 ( n2030 ) , .IN3 ( n2029 ) 
    , .IN2 ( bank_registro_registros[63] ) , .Q ( n1900 ) 
    , .IN4 ( bank_registro_registros[45] ) ) ;
AO22X1 U779 (.IN1 ( n2028 ) , .IN3 ( n2027 ) 
    , .IN2 ( bank_registro_registros[11] ) , .Q ( n1901 ) 
    , .IN4 ( bank_registro_registros[27] ) ) ;
FADDX1 U778 (.A ( coeficiente_a22_in[12] ) , .B ( in_reg_salida_v[11] ) 
    , .CI ( coeficiente_a22_in[17] ) , .CO ( DP_OP_1001J1_64_4995_n360 ) 
    , .S ( DP_OP_1001J1_64_4995_n361 ) ) ;
AO22X1 U777 (.IN1 ( n1642 ) , .IN3 ( n1640 ) 
    , .IN2 ( bank_registro_registros[64] ) , .Q ( n1904 ) 
    , .IN4 ( bank_registro_registros[46] ) ) ;
AO22X1 U776 (.IN1 ( n2028 ) , .IN3 ( n1634 ) 
    , .IN2 ( bank_registro_registros[12] ) , .Q ( n1905 ) 
    , .IN4 ( bank_registro_registros[28] ) ) ;
AO22X1 U791 (.IN1 ( n1642 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][1] ) , .Q ( n1780 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][1] ) ) ;
AO22X1 U790 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][1] ) , .Q ( n1783 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][1] ) ) ;
FADDX1 U789 (.A ( coeficiente_a22_in[14] ) , .B ( coeficiente_a22_in[7] ) 
    , .CI ( n1583 ) , .CO ( DP_OP_1001J1_64_4995_n476 ) 
    , .S ( DP_OP_1001J1_64_4995_n477 ) ) ;
INVX0 U788 (.ZN ( n1542 ) , .INP ( coeficiente_a22_in[2] ) ) ;
AO22X1 U787 (.IN1 ( n1643 ) , .IN3 ( n2029 ) 
    , .IN2 ( bank_registro_registros[53] ) , .Q ( n1932 ) 
    , .IN4 ( bank_registro_registros[35] ) ) ;
AO22X1 U786 (.IN1 ( n2028 ) , .IN3 ( n2027 ) 
    , .IN2 ( bank_registro_registros[1] ) , .Q ( n1933 ) 
    , .IN4 ( bank_registro_registros[17] ) ) ;
FADDX1 U785 (.A ( n1535 ) , .B ( DP_OP_1001J1_64_4995_n478 ) 
    , .CI ( DP_OP_1001J1_64_4995_n476 ) , .CO ( DP_OP_1001J1_64_4995_n460 ) 
    , .S ( DP_OP_1001J1_64_4995_n461 ) ) ;
INVX0 U784 (.ZN ( n1543 ) , .INP ( coeficiente_a22_in[3] ) ) ;
AO22X1 U799 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][13] ) , .Q ( n1759 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][13] ) ) ;
AO22X1 U798 (.IN1 ( n1643 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][6] ) , .Q ( n1800 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][6] ) ) ;
AO22X1 U797 (.IN1 ( n1637 ) , .IN3 ( n1634 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][6] ) , .Q ( n1801 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][6] ) ) ;
AO22X1 U796 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][4] ) , .Q ( n1792 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][4] ) ) ;
AO22X1 U795 (.IN1 ( n2028 ) , .IN3 ( n1634 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][4] ) , .Q ( n1793 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][4] ) ) ;
INVX0 U794 (.ZN ( n1533 ) , .INP ( coeficiente_a22_in[11] ) ) ;
INVX0 U793 (.ZN ( n1596 ) , .INP ( sos2_reg_entrada[8] ) ) ;
INVX0 U792 (.ZN ( n1582 ) , .INP ( sos2_reg_entrada[11] ) ) ;
INVX0 U807 (.ZN ( n1518 ) , .INP ( coeficiente_b12_H_v_out[15] ) ) ;
FADDX1 U806 (.A ( coeficiente_b12_H_v_out[14] ) , .B ( n1518 ) 
    , .CI ( DP_OP_1001J1_64_4995_n58 ) , .CO ( DP_OP_1001J1_64_4995_n54 ) 
    , .S ( DP_OP_1001J1_64_4995_n55 ) ) ;
INVX0 U805 (.ZN ( n1520 ) , .INP ( coeficiente_b12_H_v_out[16] ) ) ;
FADDX1 U804 (.A ( coeficiente_b12_H_v_out[15] ) , .B ( n1520 ) 
    , .CI ( DP_OP_1001J1_64_4995_n54 ) , .CO ( DP_OP_1001J1_64_4995_n50 ) 
    , .S ( DP_OP_1001J1_64_4995_n51 ) ) ;
INVX0 U803 (.ZN ( n1522 ) , .INP ( coeficiente_b12_H_v_out[17] ) ) ;
FADDX1 U802 (.A ( coeficiente_b12_H_v_out[16] ) , .B ( n1522 ) 
    , .CI ( DP_OP_1001J1_64_4995_n50 ) , .CO ( DP_OP_1001J1_64_4995_n46 ) 
    , .S ( DP_OP_1001J1_64_4995_n47 ) ) ;
INVX0 U801 (.ZN ( n1564 ) , .INP ( DP_OP_1002J1_65_247_n272 ) ) ;
AO22X1 U800 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][13] ) , .Q ( n1756 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][13] ) ) ;
INVX0 U815 (.ZN ( n1510 ) , .INP ( coeficiente_b12_H_v_out[11] ) ) ;
FADDX1 U814 (.A ( coeficiente_b12_H_v_out[10] ) , .B ( n1510 ) 
    , .CI ( DP_OP_1001J1_64_4995_n74 ) , .CO ( DP_OP_1001J1_64_4995_n70 ) 
    , .S ( DP_OP_1001J1_64_4995_n71 ) ) ;
INVX0 U813 (.ZN ( n1512 ) , .INP ( coeficiente_b12_H_v_out[12] ) ) ;
FADDX1 U812 (.A ( coeficiente_b12_H_v_out[11] ) , .B ( n1512 ) 
    , .CI ( DP_OP_1001J1_64_4995_n70 ) , .CO ( DP_OP_1001J1_64_4995_n66 ) 
    , .S ( DP_OP_1001J1_64_4995_n67 ) ) ;
INVX0 U811 (.ZN ( n1514 ) , .INP ( coeficiente_b12_H_v_out[13] ) ) ;
FADDX1 U810 (.A ( coeficiente_b12_H_v_out[12] ) , .B ( n1514 ) 
    , .CI ( DP_OP_1001J1_64_4995_n66 ) , .CO ( DP_OP_1001J1_64_4995_n62 ) 
    , .S ( DP_OP_1001J1_64_4995_n63 ) ) ;
INVX0 U809 (.ZN ( n1516 ) , .INP ( coeficiente_b12_H_v_out[14] ) ) ;
FADDX1 U808 (.A ( coeficiente_b12_H_v_out[13] ) , .B ( n1516 ) 
    , .CI ( DP_OP_1001J1_64_4995_n62 ) , .CO ( DP_OP_1001J1_64_4995_n58 ) 
    , .S ( DP_OP_1001J1_64_4995_n59 ) ) ;
FADDX1 U823 (.A ( coeficiente_a22_in[17] ) , .B ( partial_1[17] ) 
    , .CI ( DP_OP_1001J1_64_4995_n298 ) , .CO ( DP_OP_1001J1_64_4995_n297 ) 
    , .S ( DP_OP_1001J1_64_4995_n567 ) ) ;
INVX0 U822 (.ZN ( n1521 ) , .INP ( coeficiente_b12_L_v_out[17] ) ) ;
XOR3X1 U821 (.Q ( DP_OP_1001J1_64_4995_n568 ) , .IN2 ( partial_1[18] ) 
    , .IN1 ( coeficiente_a22_in[18] ) , .IN3 ( DP_OP_1001J1_64_4995_n297 ) ) ;
FADDX1 U820 (.A ( n1580 ) , .B ( DP_OP_1002J1_65_247_n273 ) 
    , .CI ( DP_OP_1002J1_65_247_n100 ) , .CO ( DP_OP_1002J1_65_247_n99 ) 
    , .S ( coeficiente_b12_L_v_out[17] ) ) ;
FADDX1 U819 (.A ( n1587 ) , .B ( sos2_reg_entrada[18] ) 
    , .CI ( DP_OP_1002J1_65_247_n131 ) , .CO ( DP_OP_1002J1_65_247_n127 ) 
    , .S ( DP_OP_1002J1_65_247_n130 ) ) ;
INVX0 U818 (.ZN ( n1526 ) , .INP ( coeficiente_a11_H_in[13] ) ) ;
FADDX1 U817 (.A ( n1527 ) , .B ( DP_OP_1001J1_64_4995_n126 ) 
    , .CI ( DP_OP_1001J1_64_4995_n125 ) , .CO ( DP_OP_1001J1_64_4995_n122 ) 
    , .S ( DP_OP_1001J1_64_4995_n123 ) ) ;
INVX0 U816 (.ZN ( n1508 ) , .INP ( coeficiente_b12_H_v_out[10] ) ) ;
FADDX1 U831 (.A ( coeficiente_b12_L_v_out[11] ) , .B ( n1511 ) 
    , .CI ( DP_OP_1001J1_64_4995_n217 ) , .CO ( DP_OP_1001J1_64_4995_n213 ) 
    , .S ( DP_OP_1001J1_64_4995_n214 ) ) ;
INVX0 U830 (.ZN ( n1513 ) , .INP ( coeficiente_b12_L_v_out[13] ) ) ;
FADDX1 U829 (.A ( coeficiente_a22_in[14] ) , .B ( partial_1[14] ) 
    , .CI ( DP_OP_1001J1_64_4995_n301 ) , .CO ( DP_OP_1001J1_64_4995_n300 ) 
    , .S ( DP_OP_1001J1_64_4995_n564 ) ) ;
INVX0 U828 (.ZN ( n1515 ) , .INP ( coeficiente_b12_L_v_out[14] ) ) ;
FADDX1 U827 (.A ( coeficiente_a22_in[15] ) , .B ( partial_1[15] ) 
    , .CI ( DP_OP_1001J1_64_4995_n300 ) , .CO ( DP_OP_1001J1_64_4995_n299 ) 
    , .S ( DP_OP_1001J1_64_4995_n565 ) ) ;
INVX0 U826 (.ZN ( n1517 ) , .INP ( coeficiente_b12_L_v_out[15] ) ) ;
FADDX1 U825 (.A ( coeficiente_a22_in[16] ) , .B ( partial_1[16] ) 
    , .CI ( DP_OP_1001J1_64_4995_n299 ) , .CO ( DP_OP_1001J1_64_4995_n298 ) 
    , .S ( DP_OP_1001J1_64_4995_n566 ) ) ;
INVX0 U824 (.ZN ( n1519 ) , .INP ( coeficiente_b12_L_v_out[16] ) ) ;
FADDX1 U839 (.A ( coeficiente_a22_in[1] ) , .B ( DP_OP_1001J1_64_4995_n314 ) 
    , .CI ( partial_1[1] ) , .CO ( DP_OP_1001J1_64_4995_n313 ) 
    , .S ( DP_OP_1001J1_64_4995_n551 ) ) ;
FADDX1 U838 (.A ( n1554 ) , .B ( DP_OP_1001J1_64_4995_n273 ) 
    , .CI ( DP_OP_1001J1_64_4995_n272 ) , .CO ( DP_OP_1001J1_64_4995_n269 ) 
    , .S ( DP_OP_1001J1_64_4995_n270 ) ) ;
FADDX1 U837 (.A ( coeficiente_a22_in[2] ) , .B ( DP_OP_1001J1_64_4995_n313 ) 
    , .CI ( partial_1[2] ) , .CO ( DP_OP_1001J1_64_4995_n312 ) 
    , .S ( DP_OP_1001J1_64_4995_n552 ) ) ;
FADDX1 U836 (.A ( coeficiente_a22_in[3] ) , .B ( DP_OP_1001J1_64_4995_n312 ) 
    , .CI ( partial_1[3] ) , .CO ( DP_OP_1001J1_64_4995_n311 ) 
    , .S ( DP_OP_1001J1_64_4995_n553 ) ) ;
INVX0 U835 (.ZN ( n1507 ) , .INP ( coeficiente_b12_L_v_out[10] ) ) ;
INVX0 U834 (.ZN ( n1509 ) , .INP ( coeficiente_b12_L_v_out[11] ) ) ;
FADDX1 U833 (.A ( coeficiente_b12_L_v_out[10] ) , .B ( n1509 ) 
    , .CI ( DP_OP_1001J1_64_4995_n221 ) , .CO ( DP_OP_1001J1_64_4995_n217 ) 
    , .S ( DP_OP_1001J1_64_4995_n218 ) ) ;
INVX0 U832 (.ZN ( n1511 ) , .INP ( coeficiente_b12_L_v_out[12] ) ) ;
FADDX1 U847 (.A ( n1616 ) , .B ( DP_OP_1004J1_67_3033_n37 ) 
    , .CI ( DP_OP_1004J1_67_3033_n34 ) , .CO ( DP_OP_1004J1_67_3033_n31 ) 
    , .S ( DP_OP_1004J1_67_3033_n32 ) ) ;
FADDX1 U846 (.A ( partial_3_H[18] ) , .B ( DP_OP_1004J1_67_3033_n33 ) 
    , .CI ( DP_OP_1004J1_67_3033_n30 ) , .CO ( DP_OP_1004J1_67_3033_n27 ) 
    , .S ( DP_OP_1004J1_67_3033_n28 ) ) ;
FADDX1 U845 (.A ( partial_3_H[14] ) , .B ( partial_3_H[17] ) 
    , .CI ( DP_OP_1004J1_67_3033_n29 ) , .CO ( DP_OP_1004J1_67_3033_n25 ) 
    , .S ( DP_OP_1004J1_67_3033_n26 ) ) ;
INVX0 U844 (.ZN ( n1613 ) , .INP ( partial_3_H[17] ) ) ;
INVX0 U843 (.ZN ( n1553 ) , .INP ( coeficiente_b11_L_v_out[13] ) ) ;
AO22X1 U842 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[3][0] ) , .Q ( n1740 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[2][0] ) ) ;
AO22X1 U841 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][0] ) , .Q ( n1743 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][0] ) ) ;
INVX0 U840 (.ZN ( n1559 ) , .INP ( coeficiente_b11_L_v_out[9] ) ) ;
FADDX1 U855 (.A ( partial_3_L[14] ) , .B ( partial_3_L[17] ) 
    , .CI ( DP_OP_1003J1_66_5789_n29 ) , .CO ( DP_OP_1003J1_66_5789_n25 ) 
    , .S ( DP_OP_1003J1_66_5789_n26 ) ) ;
FADDX1 U854 (.A ( partial_3_L[15] ) , .B ( n1600 ) , .CI ( partial_3_L[18] ) 
    , .CO ( DP_OP_1003J1_66_5789_n23 ) , .S ( DP_OP_1003J1_66_5789_n24 ) ) ;
INVX0 U853 (.ZN ( n1601 ) , .INP ( partial_3_L[16] ) ) ;
INVX0 U852 (.ZN ( n1600 ) , .INP ( partial_3_L[17] ) ) ;
INVX0 U851 (.ZN ( n1599 ) , .INP ( partial_3_L[18] ) ) ;
INVX0 U850 (.ZN ( n1617 ) , .INP ( partial_3_H[13] ) ) ;
INVX0 U849 (.ZN ( n1624 ) , .INP ( partial_3_H[6] ) ) ;
FADDX1 U848 (.A ( n1617 ) , .B ( DP_OP_1004J1_67_3033_n41 ) 
    , .CI ( DP_OP_1004J1_67_3033_n38 ) , .CO ( DP_OP_1004J1_67_3033_n35 ) 
    , .S ( DP_OP_1004J1_67_3033_n36 ) ) ;
AO22X1 U863 (.IN1 ( n1643 ) , .IN3 ( n1640 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][3] ) , .Q ( n1864 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][3] ) ) ;
AO22X1 U862 (.IN1 ( n1637 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][3] ) , .Q ( n1865 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][3] ) ) ;
FADDX1 U861 (.A ( n1608 ) , .B ( DP_OP_1003J1_66_5789_n61 ) 
    , .CI ( DP_OP_1003J1_66_5789_n58 ) , .CO ( DP_OP_1003J1_66_5789_n55 ) 
    , .S ( DP_OP_1003J1_66_5789_n56 ) ) ;
FADDX1 U860 (.A ( n1607 ) , .B ( DP_OP_1003J1_66_5789_n57 ) 
    , .CI ( DP_OP_1003J1_66_5789_n54 ) , .CO ( DP_OP_1003J1_66_5789_n51 ) 
    , .S ( DP_OP_1003J1_66_5789_n52 ) ) ;
FADDX1 U859 (.A ( n1606 ) , .B ( DP_OP_1003J1_66_5789_n53 ) 
    , .CI ( DP_OP_1003J1_66_5789_n50 ) , .CO ( DP_OP_1003J1_66_5789_n47 ) 
    , .S ( DP_OP_1003J1_66_5789_n48 ) ) ;
FADDX1 U858 (.A ( n1605 ) , .B ( DP_OP_1003J1_66_5789_n49 ) 
    , .CI ( DP_OP_1003J1_66_5789_n46 ) , .CO ( DP_OP_1003J1_66_5789_n43 ) 
    , .S ( DP_OP_1003J1_66_5789_n44 ) ) ;
FADDX1 U857 (.A ( n1601 ) , .B ( DP_OP_1003J1_66_5789_n37 ) 
    , .CI ( DP_OP_1003J1_66_5789_n34 ) , .CO ( DP_OP_1003J1_66_5789_n31 ) 
    , .S ( DP_OP_1003J1_66_5789_n32 ) ) ;
FADDX1 U856 (.A ( partial_3_L[18] ) , .B ( DP_OP_1003J1_66_5789_n33 ) 
    , .CI ( DP_OP_1003J1_66_5789_n30 ) , .CO ( DP_OP_1003J1_66_5789_n27 ) 
    , .S ( DP_OP_1003J1_66_5789_n28 ) ) ;
AO22X1 U871 (.IN1 ( n1642 ) , .IN3 ( n1639 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[3][10] ) , .Q ( n1968 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[2][10] ) ) ;
AO22X1 U870 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][10] ) , .Q ( n1971 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[5][10] ) ) ;
INVX0 U869 (.ZN ( n1610 ) , .INP ( partial_3_L[7] ) ) ;
AO22X1 U868 (.IN1 ( n1643 ) , .IN3 ( n1640 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[3][5] ) , .Q ( n1872 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[2][5] ) ) ;
AO22X1 U867 (.IN1 ( n1637 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][5] ) , .Q ( n1873 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][5] ) ) ;
INVX0 U866 (.ZN ( n1611 ) , .INP ( partial_3_L[6] ) ) ;
FADDX1 U865 (.A ( n1609 ) , .B ( n1611 ) , .CI ( DP_OP_1003J1_66_5789_n71 ) 
    , .CO ( DP_OP_1003J1_66_5789_n67 ) , .S ( DP_OP_1003J1_66_5789_n68 ) ) ;
INVX0 U864 (.ZN ( n1606 ) , .INP ( partial_3_L[11] ) ) ;
AND3X1 U879 (.IN2 ( seleccion_2_ ) , .IN1 ( seleccion_1_ ) , .IN3 ( n1492 ) 
    , .Q ( n2026 ) ) ;
AND3X1 U878 (.IN2 ( seleccion_1_ ) , .IN1 ( n1035 ) , .IN3 ( n1493 ) 
    , .Q ( n2029 ) ) ;
INVX0 U877 (.ZN ( n1631 ) , .INP ( n1472 ) ) ;
INVX0 U876 (.ZN ( n1642 ) , .INP ( n1645 ) ) ;
INVX0 U875 (.ZN ( n1639 ) , .INP ( n1470 ) ) ;
INVX0 U874 (.ZN ( n1632 ) , .INP ( n1472 ) ) ;
INVX0 U873 (.ZN ( n1643 ) , .INP ( n1645 ) ) ;
INVX0 U872 (.ZN ( n1640 ) , .INP ( n1470 ) ) ;
AOI22X1 U887 (.IN4 ( bank_registro_registros[139] ) 
    , .IN2 ( bank_registro_registros[103] ) , .IN3 ( n1631 ) , .IN1 ( n1627 ) 
    , .QN ( n1920 ) ) ;
FADDX1 U886 (.A ( in_reg_salida_v[15] ) , .B ( coeficiente_a22_in[16] ) 
    , .CI ( DP_OP_1001J1_64_4995_n344 ) , .CO ( DP_OP_1001J1_64_4995_n340 ) 
    , .S ( DP_OP_1001J1_64_4995_n341 ) ) ;
AO22X1 U885 (.IN1 ( n1641 ) , .IN3 ( n2029 ) 
    , .IN2 ( bank_registro_registros[68] ) , .Q ( n1921 ) 
    , .IN4 ( bank_registro_registros[50] ) ) ;
AOI22X1 U884 (.IN4 ( bank_registro_registros[140] ) 
    , .IN2 ( bank_registro_registros[104] ) , .IN3 ( n2026 ) , .IN1 ( n1626 ) 
    , .QN ( n1925 ) ) ;
FADDX1 U883 (.A ( in_reg_salida_v[16] ) , .B ( coeficiente_a22_in[17] ) 
    , .CI ( n1538 ) , .CO ( DP_OP_1001J1_64_4995_n338 ) 
    , .S ( DP_OP_1001J1_64_4995_n339 ) ) ;
AO22X1 U882 (.IN1 ( n2030 ) , .IN3 ( n2029 ) 
    , .IN2 ( bank_registro_registros[69] ) , .Q ( n1926 ) 
    , .IN4 ( bank_registro_registros[51] ) ) ;
AOI22X1 U881 (.IN4 ( bank_registro_registros[141] ) 
    , .IN2 ( bank_registro_registros[105] ) , .IN3 ( n2026 ) , .IN1 ( n1626 ) 
    , .QN ( n1930 ) ) ;
INVX0 U880 (.ZN ( n1641 ) , .INP ( n1645 ) ) ;
FADDX1 U895 (.A ( n1526 ) , .B ( DP_OP_1001J1_64_4995_n127 ) 
    , .CI ( DP_OP_1001J1_64_4995_n550 ) , .CO ( DP_OP_1001J1_64_4995_n40 ) 
    , .S ( partial_2_H[0] ) ) ;
INVX0 U894 (.ZN ( n1563 ) , .INP ( sos2_reg_entrada[0] ) ) ;
FADDX1 U893 (.A ( n1596 ) , .B ( n1582 ) , .CI ( n1533 ) 
    , .CO ( DP_OP_1001J1_64_4995_n480 ) , .S ( DP_OP_1001J1_64_4995_n481 ) ) ;
AO22X1 U892 (.IN1 ( n2030 ) , .IN3 ( n1640 ) 
    , .IN2 ( bank_registro_registros[52] ) , .Q ( n1892 ) 
    , .IN4 ( bank_registro_registros[34] ) ) ;
AO22X1 U891 (.IN1 ( n2028 ) , .IN3 ( n2027 ) 
    , .IN2 ( bank_registro_registros[0] ) , .Q ( n1893 ) 
    , .IN4 ( bank_registro_registros[16] ) ) ;
INVX0 U890 (.ZN ( n1541 ) , .INP ( coeficiente_a22_in[1] ) ) ;
FADDX1 U889 (.A ( n1540 ) , .B ( DP_OP_1001J1_64_4995_n348 ) 
    , .CI ( DP_OP_1001J1_64_4995_n345 ) , .CO ( DP_OP_1001J1_64_4995_n342 ) 
    , .S ( DP_OP_1001J1_64_4995_n343 ) ) ;
AO22X1 U888 (.IN1 ( n1644 ) , .IN3 ( n2029 ) 
    , .IN2 ( bank_registro_registros[67] ) , .Q ( n1916 ) 
    , .IN4 ( bank_registro_registros[49] ) ) ;
INVX0 U903 (.ZN ( n1612 ) , .INP ( partial_3_L[5] ) ) ;
FADDX1 U902 (.A ( n1610 ) , .B ( n1612 ) , .CI ( DP_OP_1003J1_66_5789_n72 ) 
    , .CO ( DP_OP_1003J1_66_5789_n18 ) , .S ( bajo_reg_entrada[0] ) ) ;
FADDX1 U901 (.A ( n1601 ) , .B ( DP_OP_1003J1_66_5789_n23 ) 
    , .CI ( DP_OP_1003J1_66_5789_n5 ) , .CO ( DP_OP_1003J1_66_5789_n4 ) 
    , .S ( bajo_reg_entrada[14] ) ) ;
FADDX1 U900 (.A ( partial_3_L[16] ) , .B ( n1600 ) 
    , .CI ( DP_OP_1003J1_66_5789_n4 ) , .CO ( DP_OP_1003J1_66_5789_n3 ) 
    , .S ( bajo_reg_entrada[15] ) ) ;
FADDX1 U899 (.A ( partial_3_L[17] ) , .B ( n1599 ) 
    , .CI ( DP_OP_1003J1_66_5789_n3 ) , .CO ( DP_OP_1003J1_66_5789_n2 ) 
    , .S ( bajo_reg_entrada[16] ) ) ;
INVX0 U898 (.ZN ( n1625 ) , .INP ( partial_3_H[5] ) ) ;
FADDX1 U897 (.A ( n1614 ) , .B ( DP_OP_1004J1_67_3033_n23 ) 
    , .CI ( DP_OP_1004J1_67_3033_n5 ) , .CO ( DP_OP_1004J1_67_3033_n4 ) 
    , .S ( alto_reg_entrada[14] ) ) ;
XOR3X1 U896 (.Q ( alto_reg_entrada[15] ) , .IN2 ( n1613 ) 
    , .IN1 ( partial_3_H[16] ) , .IN3 ( DP_OP_1004J1_67_3033_n4 ) ) ;
AO22X1 U911 (.IN1 ( n1641 ) , .IN3 ( n1639 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[3][15] ) , .Q ( n1988 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[2][15] ) ) ;
AO22X1 U910 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][15] ) , .Q ( n1991 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[5][15] ) ) ;
AO22X1 U909 (.IN1 ( n1641 ) , .IN3 ( n1639 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[3][16] ) , .Q ( n1992 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[2][16] ) ) ;
AO22X1 U908 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][16] ) , .Q ( n1995 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[5][16] ) ) ;
AO22X1 U907 (.IN1 ( n1642 ) , .IN3 ( n1639 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[3][17] ) , .Q ( n1996 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[2][17] ) ) ;
AO22X1 U906 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][17] ) , .Q ( n1999 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[5][17] ) ) ;
AO22X1 U905 (.IN1 ( n1641 ) , .IN3 ( n1639 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[3][18] ) , .Q ( n2000 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[2][18] ) ) ;
AO22X1 U904 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][18] ) , .Q ( n2003 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[5][18] ) ) ;
INVX2 U919 (.INP ( reset ) , .ZN ( n1663 ) ) ;
INVX2 U918 (.INP ( reset ) , .ZN ( n1661 ) ) ;
AO22X1 U917 (.IN1 ( n1642 ) , .IN3 ( n1639 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[3][13] ) , .Q ( n1980 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[2][13] ) ) ;
AO22X1 U916 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][13] ) , .Q ( n1983 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[5][13] ) ) ;
INVX2 U915 (.INP ( reset ) , .ZN ( n1660 ) ) ;
INVX2 U914 (.INP ( reset ) , .ZN ( n1662 ) ) ;
AO22X1 U913 (.IN1 ( n1642 ) , .IN3 ( n1639 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[3][14] ) , .Q ( n1984 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[2][14] ) ) ;
AO22X1 U912 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][14] ) , .Q ( n1987 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[5][14] ) ) ;
AO22X1 U927 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][8] ) , .Q ( n2023 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[5][8] ) ) ;
INVX2 U926 (.INP ( reset ) , .ZN ( n1648 ) ) ;
AO22X1 U925 (.IN1 ( n1643 ) , .IN3 ( n1640 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[3][9] ) , .Q ( n2031 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[2][9] ) ) ;
AO22X1 U924 (.IN1 ( n1637 ) , .IN3 ( n1633 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[0][9] ) , .Q ( n2032 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[1][9] ) ) ;
AO22X1 U923 (.IN1 ( n1642 ) , .IN3 ( n1639 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[3][11] ) , .Q ( n1972 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[2][11] ) ) ;
AO22X1 U922 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][11] ) , .Q ( n1975 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[5][11] ) ) ;
AO22X1 U921 (.IN1 ( n1642 ) , .IN3 ( n1639 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[3][12] ) , .Q ( n1976 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[2][12] ) ) ;
AO22X1 U920 (.IN1 ( n2024 ) , .IN3 ( n1627 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][12] ) , .Q ( n1979 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[5][12] ) ) ;
AO22X1 U935 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][4] ) , .Q ( n2007 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[5][4] ) ) ;
AO22X1 U934 (.IN1 ( n1641 ) , .IN3 ( n1639 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[3][5] ) , .Q ( n2008 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[2][5] ) ) ;
AO22X1 U933 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][5] ) , .Q ( n2011 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[5][5] ) ) ;
AO22X1 U932 (.IN1 ( n1641 ) , .IN3 ( n1639 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[3][6] ) , .Q ( n2012 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[2][6] ) ) ;
AO22X1 U931 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][6] ) , .Q ( n2015 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[5][6] ) ) ;
AO22X1 U930 (.IN1 ( n1641 ) , .IN3 ( n1639 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[3][7] ) , .Q ( n2016 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[2][7] ) ) ;
AO22X1 U929 (.IN1 ( n2024 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][7] ) , .Q ( n2019 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[5][7] ) ) ;
AO22X1 U928 (.IN1 ( n1641 ) , .IN3 ( n1639 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[3][8] ) , .Q ( n2020 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[2][8] ) ) ;
INVX0 U943 (.ZN ( n1436 ) , .INP ( seleccion_1_ ) ) ;
INVX2 U942 (.INP ( reset ) , .ZN ( n1659 ) ) ;
INVX2 U941 (.INP ( reset ) , .ZN ( n1656 ) ) ;
INVX2 U940 (.INP ( reset ) , .ZN ( n1657 ) ) ;
INVX2 U939 (.INP ( reset ) , .ZN ( n1655 ) ) ;
INVX2 U938 (.INP ( reset ) , .ZN ( n1654 ) ) ;
INVX2 U937 (.INP ( reset ) , .ZN ( n1658 ) ) ;
AO22X1 U936 (.IN1 ( n1641 ) , .IN3 ( n1639 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[3][4] ) , .Q ( n2004 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[2][4] ) ) ;
INVX0 U951 (.ZN ( n1441 ) , .INP ( seleccion_1_ ) ) ;
XOR3X1 U950 (.Q ( partial_3_H[18] ) , .IN2 ( partial_2_H[18] ) 
    , .IN1 ( coeficiente_b11_H_v_out[18] ) , .IN3 ( DP_OP_1001J1_64_4995_n3 ) ) ;
OR4X1 U949 (.IN4 ( n1440 ) , .IN2 ( n1438 ) , .Q ( sos2_reg_entrada[3] ) 
    , .IN1 ( n1437 ) , .IN3 ( n1439 ) ) ;
AO22X1 U948 (.IN1 ( \sos1_reg/bank_registro_registros[6][3] ) 
    , .IN3 ( \sos1_reg/bank_registro_registros[7][3] ) , .IN2 ( n1629 ) 
    , .Q ( n1440 ) , .IN4 ( n2026 ) ) ;
AO22X1 U947 (.IN1 ( n2024 ) , .IN3 ( \sos1_reg/bank_registro_registros[5][3] ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][3] ) , .Q ( n1439 ) 
    , .IN4 ( n1626 ) ) ;
AO22X1 U946 (.IN1 ( n1639 ) , .IN3 ( \sos1_reg/bank_registro_registros[3][3] ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[2][3] ) , .Q ( n1438 ) 
    , .IN4 ( n1641 ) ) ;
AO22X1 U945 (.IN1 ( \sos1_reg/bank_registro_registros[1][3] ) 
    , .IN3 ( \sos1_reg/bank_registro_registros[0][3] ) , .IN2 ( n1633 ) 
    , .Q ( n1437 ) , .IN4 ( n1636 ) ) ;
NAND3X0 U944 (.QN ( n1494 ) , .IN3 ( n1436 ) , .IN2 ( n1492 ) 
    , .IN1 ( seleccion_2_ ) ) ;
AND3X1 U959 (.IN2 ( n1035 ) , .IN1 ( seleccion_2_ ) , .IN3 ( n1446 ) 
    , .Q ( n2024 ) ) ;
INVX0 U958 (.ZN ( n1446 ) , .INP ( seleccion_1_ ) ) ;
OR4X1 U957 (.IN4 ( n1445 ) , .IN2 ( n1443 ) , .Q ( sos2_reg_entrada[2] ) 
    , .IN1 ( n1442 ) , .IN3 ( n1444 ) ) ;
AO22X1 U956 (.IN1 ( \sos1_reg/bank_registro_registros[6][2] ) 
    , .IN3 ( \sos1_reg/bank_registro_registros[7][2] ) , .IN2 ( n1629 ) 
    , .Q ( n1445 ) , .IN4 ( n1631 ) ) ;
AO22X1 U955 (.IN1 ( n2024 ) , .IN3 ( \sos1_reg/bank_registro_registros[5][2] ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][2] ) , .Q ( n1444 ) 
    , .IN4 ( n1626 ) ) ;
AO22X1 U954 (.IN1 ( n1639 ) , .IN3 ( \sos1_reg/bank_registro_registros[3][2] ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[2][2] ) , .Q ( n1443 ) 
    , .IN4 ( n1641 ) ) ;
AO22X1 U953 (.IN1 ( \sos1_reg/bank_registro_registros[1][2] ) 
    , .IN3 ( \sos1_reg/bank_registro_registros[0][2] ) , .IN2 ( n1633 ) 
    , .Q ( n1442 ) , .IN4 ( n1636 ) ) ;
AND3X1 U952 (.IN2 ( n1035 ) , .IN1 ( n1493 ) , .IN3 ( n1441 ) , .Q ( n2028 ) ) ;
NAND2X0 U967 (.IN1 ( n1123 ) , .IN2 ( n1122 ) 
    , .QN ( secuencia_reloj_prioridad_salida_pre_0_ ) ) ;
OR4X1 U966 (.IN4 ( n1450 ) , .IN2 ( n1448 ) , .Q ( sos2_reg_entrada[1] ) 
    , .IN1 ( n1447 ) , .IN3 ( n1449 ) ) ;
AO22X1 U965 (.IN1 ( \sos1_reg/bank_registro_registros[6][1] ) 
    , .IN3 ( \sos1_reg/bank_registro_registros[7][1] ) , .IN2 ( n1629 ) 
    , .Q ( n1450 ) , .IN4 ( n2026 ) ) ;
AO22X1 U964 (.IN1 ( n2024 ) , .IN3 ( \sos1_reg/bank_registro_registros[5][1] ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][1] ) , .Q ( n1449 ) 
    , .IN4 ( n1626 ) ) ;
AO22X1 U963 (.IN1 ( n1639 ) , .IN3 ( \sos1_reg/bank_registro_registros[3][1] ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[2][1] ) , .Q ( n1448 ) 
    , .IN4 ( n1641 ) ) ;
AO22X1 U962 (.IN1 ( \sos1_reg/bank_registro_registros[1][1] ) 
    , .IN3 ( \sos1_reg/bank_registro_registros[0][1] ) , .IN2 ( n1633 ) 
    , .Q ( n1447 ) , .IN4 ( n1636 ) ) ;
XOR3X1 U961 (.Q ( DP_OP_1001J1_64_4995_n45 ) , .IN2 ( n1496 ) 
    , .IN1 ( coeficiente_b12_H_v_out[17] ) , .IN3 ( DP_OP_1001J1_64_4995_n46 ) ) ;
XOR3X1 U960 (.Q ( n1496 ) , .IN2 ( DP_OP_1002J1_65_247_n2 ) 
    , .IN1 ( DP_OP_1002J1_65_247_n273 ) , .IN3 ( n1598 ) ) ;
AO22X1 U975 (.IN1 ( n2024 ) , .IN3 ( bank_registro_registros[105] ) 
    , .IN2 ( bank_registro_registros[87] ) , .Q ( n1455 ) , .IN4 ( n1627 ) ) ;
OR4X1 U974 (.IN4 ( n1454 ) , .IN2 ( n1452 ) , .Q ( sos2_reg_entrada[0] ) 
    , .IN1 ( n1451 ) , .IN3 ( n1453 ) ) ;
AO22X1 U973 (.IN1 ( \sos1_reg/bank_registro_registros[6][0] ) 
    , .IN3 ( \sos1_reg/bank_registro_registros[7][0] ) , .IN2 ( n2025 ) 
    , .Q ( n1454 ) , .IN4 ( n1631 ) ) ;
AO22X1 U972 (.IN1 ( n2024 ) , .IN3 ( \sos1_reg/bank_registro_registros[5][0] ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][0] ) , .Q ( n1453 ) 
    , .IN4 ( n1627 ) ) ;
AO22X1 U971 (.IN1 ( n2029 ) , .IN3 ( \sos1_reg/bank_registro_registros[3][0] ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[2][0] ) , .Q ( n1452 ) 
    , .IN4 ( n1642 ) ) ;
AO22X1 U970 (.IN1 ( \sos1_reg/bank_registro_registros[1][0] ) 
    , .IN3 ( \sos1_reg/bank_registro_registros[0][0] ) , .IN2 ( n1633 ) 
    , .Q ( n1451 ) , .IN4 ( n1636 ) ) ;
XOR3X1 U969 (.Q ( DP_OP_1001J1_64_4995_n192 ) , .IN2 ( n1495 ) 
    , .IN1 ( coeficiente_b12_L_v_out[17] ) , .IN3 ( DP_OP_1001J1_64_4995_n193 ) ) ;
INVX0 U968 (.ZN ( n1033 ) , .INP ( n1120 ) ) ;
INVX0 U983 (.ZN ( n1471 ) , .INP ( n2025 ) ) ;
INVX0 U982 (.ZN ( n1032 ) , .INP ( n1121 ) ) ;
XOR3X1 U981 (.Q ( partial_1[18] ) , .IN2 ( n1460 ) 
    , .IN1 ( DP_OP_1001J1_64_4995_n316 ) , .IN3 ( DP_OP_1001J1_64_4995_n336 ) ) ;
NOR4X0 U980 (.IN2 ( n1456 ) , .IN1 ( n1455 ) , .IN3 ( n1457 ) , .IN4 ( n1459 ) 
    , .QN ( n1460 ) ) ;
NAND2X0 U979 (.IN1 ( n1458 ) , .IN2 ( n1931 ) , .QN ( n1459 ) ) ;
NAND2X0 U978 (.IN1 ( n2029 ) , .IN2 ( bank_registro_registros[51] ) 
    , .QN ( n1458 ) ) ;
AO22X1 U977 (.IN1 ( bank_registro_registros[123] ) 
    , .IN3 ( bank_registro_registros[141] ) , .IN2 ( n2025 ) , .Q ( n1457 ) 
    , .IN4 ( n2026 ) ) ;
AO22X1 U976 (.IN1 ( bank_registro_registros[69] ) 
    , .IN3 ( bank_registro_registros[33] ) , .IN2 ( n1641 ) , .Q ( n1456 ) 
    , .IN4 ( n2027 ) ) ;
INVX2 U991 (.INP ( sos2_reg_entrada[18] ) , .ZN ( n1588 ) ) ;
INVX2 U990 (.INP ( partial_3_H[16] ) , .ZN ( n1614 ) ) ;
INVX0 U989 (.ZN ( n1635 ) , .INP ( n2027 ) ) ;
INVX2 U988 (.INP ( n1494 ) , .ZN ( n1627 ) ) ;
INVX2 U987 (.INP ( n1469 ) , .ZN ( n1628 ) ) ;
INVX0 U986 (.ZN ( n1469 ) , .INP ( n2024 ) ) ;
AND3X1 U985 (.IN2 ( n1035 ) , .IN1 ( seleccion_1_ ) , .IN3 ( seleccion_2_ ) 
    , .Q ( n2025 ) ) ;
INVX0 U984 (.ZN ( n1629 ) , .INP ( n1471 ) ) ;
INVX2 U999 (.INP ( reset ) , .ZN ( n1652 ) ) ;
INVX0 U998 (.ZN ( n1468 ) , .INP ( n2028 ) ) ;
NAND2X1 U997 (.IN2 ( bank_registro_registros[86] ) , .IN1 ( n2024 ) 
    , .QN ( n1923 ) ) ;
INVX2 U996 (.INP ( n1635 ) , .ZN ( n1634 ) ) ;
INVX2 U995 (.INP ( n1471 ) , .ZN ( n1630 ) ) ;
INVX2 U994 (.INP ( n1494 ) , .ZN ( n1626 ) ) ;
INVX0 U993 (.ZN ( n1633 ) , .INP ( n1635 ) ) ;
NAND2X1 U992 (.IN2 ( bank_registro_registros[85] ) , .IN1 ( n2024 ) 
    , .QN ( n1918 ) ) ;
OR4X1 U1007 (.IN4 ( n1984 ) , .IN2 ( n1986 ) , .Q ( sos2_reg_entrada[14] ) 
    , .IN1 ( n1987 ) , .IN3 ( n1985 ) ) ;
INVX2 U1006 (.INP ( reset ) , .ZN ( n1649 ) ) ;
INVX2 U1005 (.INP ( reset ) , .ZN ( n1647 ) ) ;
INVX2 U1004 (.INP ( reset ) , .ZN ( n1653 ) ) ;
INVX2 U1003 (.INP ( reset ) , .ZN ( n1651 ) ) ;
INVX2 U1002 (.INP ( reset ) , .ZN ( n1650 ) ) ;
NOR3X1 U1001 (.IN2 ( n1035 ) , .IN1 ( seleccion_1_ ) , .IN3 ( seleccion_2_ ) 
    , .QN ( n2027 ) ) ;
INVX2 U1000 (.INP ( reset ) , .ZN ( n1646 ) ) ;
OR4X1 U1015 (.IN4 ( n1976 ) , .IN2 ( n1978 ) , .Q ( sos2_reg_entrada[12] ) 
    , .IN1 ( n1979 ) , .IN3 ( n1977 ) ) ;
OR4X1 U1014 (.IN4 ( n1760 ) , .IN2 ( n1762 ) , .Q ( coeficiente_a22_in[14] ) 
    , .IN1 ( n1763 ) , .IN3 ( n1761 ) ) ;
OR4X1 U1013 (.IN4 ( n1776 ) , .IN2 ( n1778 ) , .Q ( coeficiente_a22_in[18] ) 
    , .IN1 ( n1779 ) , .IN3 ( n1777 ) ) ;
XOR3X1 U1012 (.Q ( partial_2_L[18] ) , .IN2 ( DP_OP_1001J1_64_4995_n568 ) 
    , .IN1 ( DP_OP_1001J1_64_4995_n192 ) , .IN3 ( DP_OP_1001J1_64_4995_n170 ) ) ;
XOR3X1 U1011 (.Q ( partial_2_H[18] ) , .IN2 ( DP_OP_1001J1_64_4995_n568 ) 
    , .IN1 ( DP_OP_1001J1_64_4995_n45 ) , .IN3 ( DP_OP_1001J1_64_4995_n23 ) ) ;
NAND2X1 U1010 (.IN2 ( bank_registro_registros[87] ) , .IN1 ( n2024 ) 
    , .QN ( n1928 ) ) ;
OR4X1 U1009 (.IN4 ( n1988 ) , .IN2 ( n1990 ) , .Q ( sos2_reg_entrada[15] ) 
    , .IN1 ( n1991 ) , .IN3 ( n1989 ) ) ;
OR4X1 U1008 (.IN4 ( n2000 ) , .IN2 ( n2002 ) , .Q ( sos2_reg_entrada[18] ) 
    , .IN1 ( n2003 ) , .IN3 ( n2001 ) ) ;
OR4X1 U1023 (.IN4 ( n1696 ) , .IN2 ( n1698 ) , .Q ( coeficiente_a11_H_in[17] ) 
    , .IN1 ( n1699 ) , .IN3 ( n1697 ) ) ;
OR4X1 U1022 (.IN4 ( n1748 ) , .IN2 ( n1750 ) , .Q ( coeficiente_a22_in[11] ) 
    , .IN1 ( n1751 ) , .IN3 ( n1749 ) ) ;
OR4X1 U1021 (.IN4 ( n1680 ) , .IN2 ( n1682 ) , .Q ( coeficiente_a11_H_in[13] ) 
    , .IN1 ( n1683 ) , .IN3 ( n1681 ) ) ;
OR4X1 U1020 (.IN4 ( n1756 ) , .IN2 ( n1758 ) , .Q ( coeficiente_a22_in[13] ) 
    , .IN1 ( n1759 ) , .IN3 ( n1757 ) ) ;
OR4X1 U1019 (.IN4 ( n1804 ) , .IN2 ( n1806 ) , .Q ( coeficiente_a22_in[7] ) 
    , .IN1 ( n1807 ) , .IN3 ( n1805 ) ) ;
OR4X1 U1018 (.IN4 ( n1832 ) , .IN2 ( n1834 ) 
    , .Q ( coeficiente_b11_L_v_out[13] ) , .IN1 ( n1835 ) , .IN3 ( n1833 ) ) ;
OR4X1 U1017 (.IN4 ( n2031 ) , .IN2 ( n2033 ) , .Q ( sos2_reg_entrada[9] ) 
    , .IN1 ( n2034 ) , .IN3 ( n2032 ) ) ;
OR4X1 U1016 (.IN4 ( n1752 ) , .IN2 ( n1754 ) , .Q ( coeficiente_a22_in[12] ) 
    , .IN1 ( n1755 ) , .IN3 ( n1753 ) ) ;
OR4X1 U1031 (.IN4 ( n1836 ) , .IN2 ( n1838 ) 
    , .Q ( coeficiente_b11_L_v_out[14] ) , .IN1 ( n1839 ) , .IN3 ( n1837 ) ) ;
OR4X1 U1030 (.IN4 ( n1772 ) , .IN2 ( n1774 ) , .Q ( coeficiente_a22_in[17] ) 
    , .IN1 ( n1775 ) , .IN3 ( n1773 ) ) ;
OR4X1 U1029 (.IN4 ( n2020 ) , .IN2 ( n2022 ) , .Q ( sos2_reg_entrada[8] ) 
    , .IN1 ( n2023 ) , .IN3 ( n2021 ) ) ;
OR4X1 U1028 (.IN4 ( n1844 ) , .IN2 ( n1846 ) 
    , .Q ( coeficiente_b11_L_v_out[16] ) , .IN1 ( n1847 ) , .IN3 ( n1845 ) ) ;
OR4X1 U1027 (.IN4 ( n1812 ) , .IN2 ( n1814 ) , .Q ( coeficiente_a22_in[9] ) 
    , .IN1 ( n1815 ) , .IN3 ( n1813 ) ) ;
OR4X1 U1026 (.IN4 ( n1744 ) , .IN2 ( n1746 ) , .Q ( coeficiente_a22_in[10] ) 
    , .IN1 ( n1747 ) , .IN3 ( n1745 ) ) ;
OR4X1 U1025 (.IN4 ( n1768 ) , .IN2 ( n1770 ) , .Q ( coeficiente_a22_in[16] ) 
    , .IN1 ( n1771 ) , .IN3 ( n1769 ) ) ;
OR4X1 U1024 (.IN4 ( n1840 ) , .IN2 ( n1842 ) 
    , .Q ( coeficiente_b11_L_v_out[15] ) , .IN1 ( n1843 ) , .IN3 ( n1841 ) ) ;
NAND2X1 U1039 (.IN2 ( bank_registro_registros[15] ) , .IN1 ( n1638 ) 
    , .QN ( n1931 ) ) ;
OR4X1 U1038 (.IN4 ( n1764 ) , .IN2 ( n1766 ) , .Q ( coeficiente_a22_in[15] ) 
    , .IN1 ( n1767 ) , .IN3 ( n1765 ) ) ;
OR4X1 U1037 (.IN4 ( n1972 ) , .IN2 ( n1974 ) , .Q ( sos2_reg_entrada[11] ) 
    , .IN1 ( n1975 ) , .IN3 ( n1973 ) ) ;
OR4X1 U1036 (.IN4 ( n1800 ) , .IN2 ( n1802 ) , .Q ( coeficiente_a22_in[6] ) 
    , .IN1 ( n1803 ) , .IN3 ( n1801 ) ) ;
OR4X1 U1035 (.IN4 ( n1684 ) , .IN2 ( n1686 ) , .Q ( coeficiente_a11_H_in[14] ) 
    , .IN1 ( n1687 ) , .IN3 ( n1685 ) ) ;
OR4X1 U1034 (.IN4 ( n1848 ) , .IN2 ( n1850 ) 
    , .Q ( coeficiente_b11_L_v_out[17] ) , .IN1 ( n1851 ) , .IN3 ( n1849 ) ) ;
OR4X1 U1033 (.IN4 ( n1980 ) , .IN2 ( n1982 ) , .Q ( sos2_reg_entrada[13] ) 
    , .IN1 ( n1983 ) , .IN3 ( n1981 ) ) ;
OR4X1 U1032 (.IN4 ( n1968 ) , .IN2 ( n1970 ) , .Q ( sos2_reg_entrada[10] ) 
    , .IN1 ( n1971 ) , .IN3 ( n1969 ) ) ;
INVX0 U1047 (.ZN ( n1637 ) , .INP ( n1468 ) ) ;
INVX0 U1046 (.ZN ( n1636 ) , .INP ( n1468 ) ) ;
INVX0 U1045 (.ZN ( n1638 ) , .INP ( n1468 ) ) ;
NOR3X0 U1044 (.IN2 ( seleccion_2_ ) , .QN ( n2030 ) , .IN1 ( n1035 ) 
    , .IN3 ( n1491 ) ) ;
INVX0 U1043 (.ZN ( n1645 ) , .INP ( n2030 ) ) ;
OR4X1 U1042 (.IN4 ( n1996 ) , .IN2 ( n1998 ) , .Q ( sos2_reg_entrada[17] ) 
    , .IN1 ( n1999 ) , .IN3 ( n1997 ) ) ;
INVX2 U1041 (.INP ( sos2_reg_entrada[17] ) , .ZN ( n1587 ) ) ;
OR4X1 U1040 (.IN4 ( n1992 ) , .IN2 ( n1994 ) , .Q ( sos2_reg_entrada[16] ) 
    , .IN1 ( n1995 ) , .IN3 ( n1993 ) ) ;
AO22X1 U1055 (.IN1 ( n1636 ) , .IN3 ( n1633 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[0][18] ) , .Q ( n2001 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[1][18] ) ) ;
AO22X1 U1054 (.IN1 ( n1636 ) , .IN3 ( n1633 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[0][16] ) , .Q ( n1993 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[1][16] ) ) ;
OR4X1 U1053 (.IN4 ( n2016 ) , .IN2 ( n2018 ) , .Q ( sos2_reg_entrada[7] ) 
    , .IN1 ( n2019 ) , .IN3 ( n2017 ) ) ;
OR4X1 U1052 (.IN4 ( n2012 ) , .IN2 ( n2014 ) , .Q ( sos2_reg_entrada[6] ) 
    , .IN1 ( n2015 ) , .IN3 ( n2013 ) ) ;
OR4X1 U1051 (.IN4 ( n2008 ) , .IN2 ( n2010 ) , .Q ( sos2_reg_entrada[5] ) 
    , .IN1 ( n2011 ) , .IN3 ( n2009 ) ) ;
OR4X1 U1050 (.IN4 ( n2004 ) , .IN2 ( n2006 ) , .Q ( sos2_reg_entrada[4] ) 
    , .IN1 ( n2007 ) , .IN3 ( n2005 ) ) ;
AND2X1 U1049 (.IN1 ( n1526 ) , .IN2 ( n1489 ) , .Q ( n1476 ) ) ;
INVX0 U1048 (.ZN ( bajo_reg_entrada[18] ) , .INP ( DP_OP_1003J1_66_5789_n2 ) ) ;
AND2X1 U1063 (.IN1 ( n1498 ) , .IN2 ( n1480 ) , .Q ( n1481 ) ) ;
AND2X1 U1062 (.IN1 ( n1497 ) , .IN2 ( n1479 ) , .Q ( n1480 ) ) ;
AND2X1 U1061 (.IN1 ( n1505 ) , .IN2 ( n1478 ) , .Q ( n1479 ) ) ;
AND2X1 U1060 (.IN1 ( n1504 ) , .IN2 ( n1477 ) , .Q ( n1478 ) ) ;
AND2X1 U1059 (.IN1 ( n1503 ) , .IN2 ( n1506 ) , .Q ( n1477 ) ) ;
AND2X1 U1058 (.IN1 ( n1528 ) , .IN2 ( n1485 ) , .Q ( n1475 ) ) ;
AND2X1 U1057 (.IN1 ( n1502 ) , .IN2 ( n1484 ) , .Q ( n1474 ) ) ;
AO22X1 U1056 (.IN1 ( n1636 ) , .IN3 ( n1633 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[0][17] ) , .Q ( n1997 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[1][17] ) ) ;
AND2X1 U1071 (.IN1 ( n1525 ) , .IN2 ( n1488 ) , .Q ( n1489 ) ) ;
AND2X1 U1070 (.IN1 ( n1524 ) , .IN2 ( n1487 ) , .Q ( n1488 ) ) ;
AND2X1 U1069 (.IN1 ( n1523 ) , .IN2 ( n1474 ) , .Q ( n1487 ) ) ;
AND2X1 U1068 (.IN1 ( n1529 ) , .IN2 ( n1475 ) , .Q ( n1486 ) ) ;
AND2X1 U1067 (.IN1 ( n1527 ) , .IN2 ( n1476 ) , .Q ( n1485 ) ) ;
AND2X1 U1066 (.IN1 ( n1501 ) , .IN2 ( n1483 ) , .Q ( n1484 ) ) ;
AND2X1 U1065 (.IN1 ( n1500 ) , .IN2 ( n1482 ) , .Q ( n1483 ) ) ;
AND2X1 U1064 (.IN1 ( n1499 ) , .IN2 ( n1481 ) , .Q ( n1482 ) ) ;
NOR4X0 U1079 (.IN2 ( n1738 ) , .IN1 ( n1739 ) , .IN3 ( n1737 ) , .IN4 ( n1736 ) 
    , .QN ( n1502 ) ) ;
NOR4X0 U1078 (.IN2 ( n1734 ) , .IN1 ( n1735 ) , .IN3 ( n1733 ) , .IN4 ( n1732 ) 
    , .QN ( n1501 ) ) ;
NOR4X0 U1077 (.IN2 ( n1730 ) , .IN1 ( n1731 ) , .IN3 ( n1729 ) , .IN4 ( n1728 ) 
    , .QN ( n1500 ) ) ;
NOR4X0 U1076 (.IN2 ( n1726 ) , .IN1 ( n1727 ) , .IN3 ( n1725 ) , .IN4 ( n1724 ) 
    , .QN ( n1499 ) ) ;
NOR4X0 U1075 (.IN2 ( n1722 ) , .IN1 ( n1723 ) , .IN3 ( n1721 ) , .IN4 ( n1720 ) 
    , .QN ( n1498 ) ) ;
NOR4X0 U1074 (.IN2 ( n1718 ) , .IN1 ( n1719 ) , .IN3 ( n1717 ) , .IN4 ( n1716 ) 
    , .QN ( n1497 ) ) ;
XOR3X1 U1073 (.Q ( n1495 ) , .IN2 ( DP_OP_1002J1_65_247_n127 ) 
    , .IN1 ( DP_OP_1002J1_65_247_n99 ) , .IN3 ( n1598 ) ) ;
AND2X1 U1072 (.IN1 ( n1530 ) , .IN2 ( n1486 ) , .Q ( n1490 ) ) ;
XOR2X1 U1087 (.IN2 ( n1480 ) , .Q ( coeficiente_b11_H_v_out[5] ) 
    , .IN1 ( n1498 ) ) ;
XOR2X1 U1086 (.IN2 ( n1479 ) , .Q ( coeficiente_b11_H_v_out[4] ) 
    , .IN1 ( n1497 ) ) ;
XOR2X1 U1085 (.IN2 ( n1478 ) , .Q ( coeficiente_b11_H_v_out[3] ) 
    , .IN1 ( n1505 ) ) ;
XOR2X1 U1084 (.IN2 ( n1477 ) , .Q ( coeficiente_b11_H_v_out[2] ) 
    , .IN1 ( n1504 ) ) ;
XOR2X1 U1083 (.IN2 ( n1506 ) , .Q ( coeficiente_b11_H_v_out[1] ) 
    , .IN1 ( n1503 ) ) ;
NOR4X0 U1082 (.IN2 ( n1714 ) , .IN1 ( n1715 ) , .IN3 ( n1713 ) , .IN4 ( n1712 ) 
    , .QN ( n1505 ) ) ;
NOR4X0 U1081 (.IN2 ( n1710 ) , .IN1 ( n1711 ) , .IN3 ( n1709 ) , .IN4 ( n1708 ) 
    , .QN ( n1504 ) ) ;
NOR4X0 U1080 (.IN2 ( n1706 ) , .IN1 ( n1707 ) , .IN3 ( n1705 ) , .IN4 ( n1704 ) 
    , .QN ( n1503 ) ) ;
XOR2X1 U1095 (.IN2 ( n1489 ) , .Q ( coeficiente_b11_H_v_out[13] ) 
    , .IN1 ( n1526 ) ) ;
XOR2X1 U1094 (.IN2 ( n1488 ) , .Q ( coeficiente_b11_H_v_out[12] ) 
    , .IN1 ( n1525 ) ) ;
XOR2X1 U1093 (.IN2 ( n1487 ) , .Q ( coeficiente_b11_H_v_out[11] ) 
    , .IN1 ( n1524 ) ) ;
XOR2X1 U1092 (.IN2 ( n1474 ) , .Q ( coeficiente_b11_H_v_out[10] ) 
    , .IN1 ( n1523 ) ) ;
XOR2X1 U1091 (.IN2 ( n1484 ) , .Q ( coeficiente_b11_H_v_out[9] ) 
    , .IN1 ( n1502 ) ) ;
XOR2X1 U1090 (.IN2 ( n1483 ) , .Q ( coeficiente_b11_H_v_out[8] ) 
    , .IN1 ( n1501 ) ) ;
XOR2X1 U1089 (.IN2 ( n1482 ) , .Q ( coeficiente_b11_H_v_out[7] ) 
    , .IN1 ( n1500 ) ) ;
XOR2X1 U1088 (.IN2 ( n1481 ) , .Q ( coeficiente_b11_H_v_out[6] ) 
    , .IN1 ( n1499 ) ) ;
AO222X1 U1103 (.Q ( DP_OP_1001J1_64_4995_n166 ) 
    , .IN2 ( coeficiente_b11_L_v_out[1] ) , .IN1 ( n1561 ) , .IN3 ( n1561 ) 
    , .IN4 ( partial_2_L[1] ) , .IN6 ( partial_2_L[1] ) 
    , .IN5 ( coeficiente_b11_L_v_out[1] ) ) ;
AND2X1 U1102 (.IN1 ( partial_2_H[0] ) , .IN2 ( coeficiente_b11_H_v_out[0] ) 
    , .Q ( n1562 ) ) ;
AND2X1 U1101 (.IN1 ( partial_2_L[0] ) , .IN2 ( coeficiente_b11_L_v_out[0] ) 
    , .Q ( n1561 ) ) ;
XOR2X1 U1100 (.IN2 ( n1490 ) , .Q ( coeficiente_b11_H_v_out[18] ) 
    , .IN1 ( n1531 ) ) ;
XOR2X1 U1099 (.IN2 ( n1486 ) , .Q ( coeficiente_b11_H_v_out[17] ) 
    , .IN1 ( n1530 ) ) ;
XOR2X1 U1098 (.IN2 ( n1475 ) , .Q ( coeficiente_b11_H_v_out[16] ) 
    , .IN1 ( n1529 ) ) ;
XOR2X1 U1097 (.IN2 ( n1485 ) , .Q ( coeficiente_b11_H_v_out[15] ) 
    , .IN1 ( n1528 ) ) ;
XOR2X1 U1096 (.IN2 ( n1476 ) , .Q ( coeficiente_b11_H_v_out[14] ) 
    , .IN1 ( n1527 ) ) ;
OR2X1 U1111 (.IN2 ( n1621 ) , .IN1 ( partial_3_H[4] ) 
    , .Q ( DP_OP_1004J1_67_3033_n77 ) ) ;
MUX21X1 U1110 (.S ( partial_3_H[4] ) , .IN2 ( n1621 ) , .IN1 ( partial_3_H[9] ) 
    , .Q ( DP_OP_1004J1_67_3033_n78 ) ) ;
OR2X1 U1109 (.IN2 ( partial_3_L[3] ) , .IN1 ( partial_3_L[11] ) 
    , .Q ( DP_OP_1003J1_66_5789_n69 ) ) ;
MUX21X1 U1108 (.S ( partial_3_L[3] ) , .IN2 ( partial_3_L[11] ) 
    , .IN1 ( n1606 ) , .Q ( DP_OP_1003J1_66_5789_n70 ) ) ;
XNOR3X1 U1107 (.Q ( n1598 ) , .IN3 ( DP_OP_1002J1_65_247_n182 ) 
    , .IN2 ( DP_OP_1002J1_65_247_n163 ) , .IN1 ( sos2_reg_entrada[17] ) ) ;
OR2X1 U1106 (.IN2 ( in_reg_salida_v[2] ) , .IN1 ( coeficiente_a22_in[15] ) 
    , .Q ( DP_OP_1001J1_64_4995_n466 ) ) ;
MUX21X1 U1105 (.S ( in_reg_salida_v[2] ) , .IN2 ( coeficiente_a22_in[15] ) 
    , .IN1 ( n1537 ) , .Q ( DP_OP_1001J1_64_4995_n467 ) ) ;
AO222X1 U1104 (.Q ( DP_OP_1001J1_64_4995_n19 ) 
    , .IN2 ( coeficiente_b11_H_v_out[1] ) , .IN1 ( n1562 ) , .IN3 ( n1562 ) 
    , .IN4 ( partial_2_H[1] ) , .IN6 ( partial_2_H[1] ) 
    , .IN5 ( coeficiente_b11_H_v_out[1] ) ) ;
AO22X1 U1119 (.IN1 ( n1638 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][11] ) , .Q ( n1673 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][11] ) ) ;
AO22X1 U1118 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][11] ) , .Q ( n1674 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][11] ) ) ;
OR4X1 U1117 (.IN4 ( n1668 ) , .IN2 ( n1670 ) , .Q ( coeficiente_a11_H_in[10] ) 
    , .IN1 ( n1671 ) , .IN3 ( n1669 ) ) ;
AO22X1 U1116 (.IN1 ( n1638 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][10] ) , .Q ( n1669 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][10] ) ) ;
AO22X1 U1115 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][10] ) , .Q ( n1670 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][10] ) ) ;
OR4X1 U1114 (.IN4 ( n1664 ) , .IN2 ( n1666 ) 
    , .Q ( coeficiente_b11_H_v_out[0] ) , .IN1 ( n1667 ) , .IN3 ( n1665 ) ) ;
AO22X1 U1113 (.IN1 ( n1636 ) , .IN3 ( n1633 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][0] ) , .Q ( n1665 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][0] ) ) ;
AO22X1 U1112 (.IN1 ( n2026 ) , .IN3 ( n1629 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][0] ) , .Q ( n1666 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][0] ) ) ;
AO22X1 U1127 (.IN1 ( n1638 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][14] ) , .Q ( n1685 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][14] ) ) ;
AO22X1 U1126 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][14] ) , .Q ( n1686 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][14] ) ) ;
AO22X1 U1125 (.IN1 ( n1638 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][13] ) , .Q ( n1681 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][13] ) ) ;
AO22X1 U1124 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][13] ) , .Q ( n1682 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][13] ) ) ;
OR4X1 U1123 (.IN4 ( n1676 ) , .IN2 ( n1678 ) , .Q ( coeficiente_a11_H_in[12] ) 
    , .IN1 ( n1679 ) , .IN3 ( n1677 ) ) ;
AO22X1 U1122 (.IN1 ( n1638 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][12] ) , .Q ( n1677 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][12] ) ) ;
AO22X1 U1121 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][12] ) , .Q ( n1678 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][12] ) ) ;
OR4X1 U1120 (.IN4 ( n1672 ) , .IN2 ( n1674 ) , .Q ( coeficiente_a11_H_in[11] ) 
    , .IN1 ( n1675 ) , .IN3 ( n1673 ) ) ;
AO22X1 U1135 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][17] ) , .Q ( n1697 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][17] ) ) ;
AO22X1 U1134 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][17] ) , .Q ( n1698 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][17] ) ) ;
OR4X1 U1133 (.IN4 ( n1692 ) , .IN2 ( n1694 ) , .Q ( coeficiente_a11_H_in[16] ) 
    , .IN1 ( n1695 ) , .IN3 ( n1693 ) ) ;
AO22X1 U1132 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][16] ) , .Q ( n1693 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][16] ) ) ;
AO22X1 U1131 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][16] ) , .Q ( n1694 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][16] ) ) ;
OR4X1 U1130 (.IN4 ( n1688 ) , .IN2 ( n1690 ) , .Q ( coeficiente_a11_H_in[15] ) 
    , .IN1 ( n1691 ) , .IN3 ( n1689 ) ) ;
AO22X1 U1129 (.IN1 ( n1638 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][15] ) , .Q ( n1689 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][15] ) ) ;
AO22X1 U1128 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][15] ) , .Q ( n1690 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][15] ) ) ;
AO22X1 U1143 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][3] ) , .Q ( n1714 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][3] ) ) ;
AO22X1 U1142 (.IN1 ( n1638 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][2] ) , .Q ( n1709 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][2] ) ) ;
AO22X1 U1141 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][2] ) , .Q ( n1710 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][2] ) ) ;
AO22X1 U1140 (.IN1 ( n1638 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][1] ) , .Q ( n1705 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][1] ) ) ;
AO22X1 U1139 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][1] ) , .Q ( n1706 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][1] ) ) ;
OR4X1 U1138 (.IN4 ( n1700 ) , .IN2 ( n1702 ) , .Q ( coeficiente_a11_H_in[18] ) 
    , .IN1 ( n1703 ) , .IN3 ( n1701 ) ) ;
AO22X1 U1137 (.IN1 ( n1638 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][18] ) , .Q ( n1701 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][18] ) ) ;
AO22X1 U1136 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][18] ) , .Q ( n1702 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][18] ) ) ;
AO22X1 U1151 (.IN1 ( n2026 ) , .IN3 ( n1629 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][7] ) , .Q ( n1730 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][7] ) ) ;
AO22X1 U1150 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][6] ) , .Q ( n1725 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][6] ) ) ;
AO22X1 U1149 (.IN1 ( n2026 ) , .IN3 ( n1629 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][6] ) , .Q ( n1726 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][6] ) ) ;
AO22X1 U1148 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][5] ) , .Q ( n1721 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][5] ) ) ;
AO22X1 U1147 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][5] ) , .Q ( n1722 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][5] ) ) ;
AO22X1 U1146 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][4] ) , .Q ( n1717 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][4] ) ) ;
AO22X1 U1145 (.IN1 ( n2026 ) , .IN3 ( n1629 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][4] ) , .Q ( n1718 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][4] ) ) ;
AO22X1 U1144 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][3] ) , .Q ( n1713 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][3] ) ) ;
OR4X1 U1159 (.IN4 ( n1740 ) , .IN2 ( n1742 ) , .Q ( coeficiente_a22_in[0] ) 
    , .IN1 ( n1743 ) , .IN3 ( n1741 ) ) ;
AO22X1 U1158 (.IN1 ( n1638 ) , .IN3 ( n2027 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][0] ) , .Q ( n1741 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][0] ) ) ;
AO22X1 U1157 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][0] ) , .Q ( n1742 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][0] ) ) ;
AO22X1 U1156 (.IN1 ( n1638 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][9] ) , .Q ( n1737 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][9] ) ) ;
AO22X1 U1155 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][9] ) , .Q ( n1738 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][9] ) ) ;
AO22X1 U1154 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][8] ) , .Q ( n1733 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][8] ) ) ;
AO22X1 U1153 (.IN1 ( n2026 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[7][8] ) , .Q ( n1734 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[6][8] ) ) ;
AO22X1 U1152 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \pos_H_reg/bank_registro_registros[0][7] ) , .Q ( n1729 ) 
    , .IN4 ( \pos_H_reg/bank_registro_registros[1][7] ) ) ;
AO22X1 U1167 (.IN1 ( n1638 ) , .IN3 ( n2027 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][13] ) , .Q ( n1757 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][13] ) ) ;
AO22X1 U1166 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][13] ) , .Q ( n1758 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][13] ) ) ;
AO22X1 U1165 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][12] ) , .Q ( n1753 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][12] ) ) ;
AO22X1 U1164 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][12] ) , .Q ( n1754 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][12] ) ) ;
AO22X1 U1163 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][11] ) , .Q ( n1749 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][11] ) ) ;
AO22X1 U1162 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][11] ) , .Q ( n1750 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][11] ) ) ;
AO22X1 U1161 (.IN1 ( n1638 ) , .IN3 ( n2027 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][10] ) , .Q ( n1745 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][10] ) ) ;
AO22X1 U1160 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][10] ) , .Q ( n1746 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][10] ) ) ;
AO22X1 U1175 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][17] ) , .Q ( n1773 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][17] ) ) ;
AO22X1 U1174 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][17] ) , .Q ( n1774 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][17] ) ) ;
AO22X1 U1173 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][16] ) , .Q ( n1769 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][16] ) ) ;
AO22X1 U1172 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][16] ) , .Q ( n1770 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][16] ) ) ;
AO22X1 U1171 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][15] ) , .Q ( n1765 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][15] ) ) ;
AO22X1 U1170 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][15] ) , .Q ( n1766 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][15] ) ) ;
AO22X1 U1169 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][14] ) , .Q ( n1761 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][14] ) ) ;
AO22X1 U1168 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][14] ) , .Q ( n1762 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][14] ) ) ;
OR4X1 U1183 (.IN4 ( n1784 ) , .IN2 ( n1786 ) , .Q ( coeficiente_a22_in[2] ) 
    , .IN1 ( n1787 ) , .IN3 ( n1785 ) ) ;
AO22X1 U1182 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][2] ) , .Q ( n1785 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][2] ) ) ;
AO22X1 U1181 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][2] ) , .Q ( n1786 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][2] ) ) ;
OR4X1 U1180 (.IN4 ( n1780 ) , .IN2 ( n1782 ) , .Q ( coeficiente_a22_in[1] ) 
    , .IN1 ( n1783 ) , .IN3 ( n1781 ) ) ;
AO22X1 U1179 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][1] ) , .Q ( n1781 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][1] ) ) ;
AO22X1 U1178 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][1] ) , .Q ( n1782 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][1] ) ) ;
AO22X1 U1177 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][18] ) , .Q ( n1777 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][18] ) ) ;
AO22X1 U1176 (.IN1 ( n2026 ) , .IN3 ( n1630 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][18] ) , .Q ( n1778 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][18] ) ) ;
AO22X1 U1191 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][5] ) , .Q ( n1798 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][5] ) ) ;
AO22X1 U1190 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][5] ) , .Q ( n1799 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][5] ) ) ;
OR4X1 U1189 (.IN4 ( n1792 ) , .IN2 ( n1794 ) , .Q ( coeficiente_a22_in[4] ) 
    , .IN1 ( n1795 ) , .IN3 ( n1793 ) ) ;
AO22X1 U1188 (.IN1 ( n1632 ) , .IN3 ( n1630 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][4] ) , .Q ( n1794 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][4] ) ) ;
AO22X1 U1187 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][4] ) , .Q ( n1795 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][4] ) ) ;
OR4X1 U1186 (.IN4 ( n1788 ) , .IN2 ( n1790 ) , .Q ( coeficiente_a22_in[3] ) 
    , .IN1 ( n1791 ) , .IN3 ( n1789 ) ) ;
AO22X1 U1185 (.IN1 ( n1638 ) , .IN3 ( n1634 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[0][3] ) , .Q ( n1789 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[1][3] ) ) ;
AO22X1 U1184 (.IN1 ( n1632 ) , .IN3 ( n1630 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][3] ) , .Q ( n1790 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][3] ) ) ;
OR4X1 U1199 (.IN4 ( n1808 ) , .IN2 ( n1810 ) , .Q ( coeficiente_a22_in[8] ) 
    , .IN1 ( n1811 ) , .IN3 ( n1809 ) ) ;
AO22X1 U1198 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][8] ) , .Q ( n1810 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][8] ) ) ;
AO22X1 U1197 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][8] ) , .Q ( n1811 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][8] ) ) ;
AO22X1 U1196 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][7] ) , .Q ( n1806 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][7] ) ) ;
AO22X1 U1195 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][7] ) , .Q ( n1807 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][7] ) ) ;
AO22X1 U1194 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][6] ) , .Q ( n1802 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][6] ) ) ;
AO22X1 U1193 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][6] ) , .Q ( n1803 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][6] ) ) ;
OR4X1 U1192 (.IN4 ( n1796 ) , .IN2 ( n1798 ) , .Q ( coeficiente_a22_in[5] ) 
    , .IN1 ( n1799 ) , .IN3 ( n1797 ) ) ;
OR4X1 U1207 (.IN4 ( n1820 ) , .IN2 ( n1822 ) 
    , .Q ( coeficiente_b11_L_v_out[10] ) , .IN1 ( n1823 ) , .IN3 ( n1821 ) ) ;
AO22X1 U1206 (.IN1 ( n2026 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][10] ) , .Q ( n1822 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][10] ) ) ;
AO22X1 U1205 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][10] ) , .Q ( n1823 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][10] ) ) ;
OR4X1 U1204 (.IN4 ( n1816 ) , .IN2 ( n1818 ) 
    , .Q ( coeficiente_b11_L_v_out[0] ) , .IN1 ( n1819 ) , .IN3 ( n1817 ) ) ;
AO22X1 U1203 (.IN1 ( n2026 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][0] ) , .Q ( n1818 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][0] ) ) ;
AO22X1 U1202 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][0] ) , .Q ( n1819 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][0] ) ) ;
AO22X1 U1201 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[7][9] ) , .Q ( n1814 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[6][9] ) ) ;
AO22X1 U1200 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos2_reg/bank_registro_registros[4][9] ) , .Q ( n1815 ) 
    , .IN4 ( \sos2_reg/bank_registro_registros[5][9] ) ) ;
AO22X1 U1215 (.IN1 ( n2026 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][13] ) , .Q ( n1834 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][13] ) ) ;
AO22X1 U1214 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][13] ) , .Q ( n1835 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][13] ) ) ;
OR4X1 U1213 (.IN4 ( n1828 ) , .IN2 ( n1830 ) 
    , .Q ( coeficiente_b11_L_v_out[12] ) , .IN1 ( n1831 ) , .IN3 ( n1829 ) ) ;
AO22X1 U1212 (.IN1 ( n2026 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][12] ) , .Q ( n1830 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][12] ) ) ;
AO22X1 U1211 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][12] ) , .Q ( n1831 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][12] ) ) ;
OR4X1 U1210 (.IN4 ( n1824 ) , .IN2 ( n1826 ) 
    , .Q ( coeficiente_b11_L_v_out[11] ) , .IN1 ( n1827 ) , .IN3 ( n1825 ) ) ;
AO22X1 U1209 (.IN1 ( n2026 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][11] ) , .Q ( n1826 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][11] ) ) ;
AO22X1 U1208 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][11] ) , .Q ( n1827 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][11] ) ) ;
AO22X1 U1223 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][17] ) , .Q ( n1851 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][17] ) ) ;
AO22X1 U1222 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][16] ) , .Q ( n1846 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][16] ) ) ;
AO22X1 U1221 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][16] ) , .Q ( n1847 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][16] ) ) ;
AO22X1 U1220 (.IN1 ( n1637 ) , .IN3 ( n2027 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[0][15] ) , .Q ( n1841 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[1][15] ) ) ;
AO22X1 U1219 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][15] ) , .Q ( n1842 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][15] ) ) ;
AO22X1 U1218 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][15] ) , .Q ( n1843 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][15] ) ) ;
AO22X1 U1217 (.IN1 ( n2026 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][14] ) , .Q ( n1838 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][14] ) ) ;
AO22X1 U1216 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][14] ) , .Q ( n1839 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][14] ) ) ;
AO22X1 U1231 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][2] ) , .Q ( n1863 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][2] ) ) ;
OR4X1 U1230 (.IN4 ( n1856 ) , .IN2 ( n1858 ) 
    , .Q ( coeficiente_b11_L_v_out[1] ) , .IN1 ( n1859 ) , .IN3 ( n1857 ) ) ;
AO22X1 U1229 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][1] ) , .Q ( n1858 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][1] ) ) ;
AO22X1 U1228 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][1] ) , .Q ( n1859 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][1] ) ) ;
OR4X1 U1227 (.IN4 ( n1852 ) , .IN2 ( n1854 ) 
    , .Q ( coeficiente_b11_L_v_out[18] ) , .IN1 ( n1855 ) , .IN3 ( n1853 ) ) ;
AO22X1 U1226 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][18] ) , .Q ( n1854 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][18] ) ) ;
AO22X1 U1225 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][18] ) , .Q ( n1855 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][18] ) ) ;
AO22X1 U1224 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][17] ) , .Q ( n1850 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][17] ) ) ;
OR4X1 U1239 (.IN4 ( n1868 ) , .IN2 ( n1870 ) 
    , .Q ( coeficiente_b11_L_v_out[4] ) , .IN1 ( n1871 ) , .IN3 ( n1869 ) ) ;
AO22X1 U1238 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][4] ) , .Q ( n1870 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][4] ) ) ;
AO22X1 U1237 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][4] ) , .Q ( n1871 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][4] ) ) ;
OR4X1 U1236 (.IN4 ( n1864 ) , .IN2 ( n1866 ) 
    , .Q ( coeficiente_b11_L_v_out[3] ) , .IN1 ( n1867 ) , .IN3 ( n1865 ) ) ;
AO22X1 U1235 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][3] ) , .Q ( n1866 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][3] ) ) ;
AO22X1 U1234 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][3] ) , .Q ( n1867 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][3] ) ) ;
OR4X1 U1233 (.IN4 ( n1860 ) , .IN2 ( n1862 ) 
    , .Q ( coeficiente_b11_L_v_out[2] ) , .IN1 ( n1863 ) , .IN3 ( n1861 ) ) ;
AO22X1 U1232 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][2] ) , .Q ( n1862 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][2] ) ) ;
AO22X1 U1247 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][7] ) , .Q ( n1882 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][7] ) ) ;
AO22X1 U1246 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][7] ) , .Q ( n1883 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][7] ) ) ;
OR4X1 U1245 (.IN4 ( n1876 ) , .IN2 ( n1878 ) 
    , .Q ( coeficiente_b11_L_v_out[6] ) , .IN1 ( n1879 ) , .IN3 ( n1877 ) ) ;
AO22X1 U1244 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][6] ) , .Q ( n1878 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][6] ) ) ;
AO22X1 U1243 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][6] ) , .Q ( n1879 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][6] ) ) ;
OR4X1 U1242 (.IN4 ( n1872 ) , .IN2 ( n1874 ) 
    , .Q ( coeficiente_b11_L_v_out[5] ) , .IN1 ( n1875 ) , .IN3 ( n1873 ) ) ;
AO22X1 U1241 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][5] ) , .Q ( n1874 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][5] ) ) ;
AO22X1 U1240 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][5] ) , .Q ( n1875 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][5] ) ) ;
AO22X1 U1255 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( bank_registro_registros[70] ) , .Q ( n1895 ) 
    , .IN4 ( bank_registro_registros[88] ) ) ;
OR4X1 U1254 (.IN4 ( n1888 ) , .IN2 ( n1890 ) 
    , .Q ( coeficiente_b11_L_v_out[9] ) , .IN1 ( n1891 ) , .IN3 ( n1889 ) ) ;
AO22X1 U1253 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][9] ) , .Q ( n1890 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][9] ) ) ;
AO22X1 U1252 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][9] ) , .Q ( n1891 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][9] ) ) ;
OR4X1 U1251 (.IN4 ( n1884 ) , .IN2 ( n1886 ) 
    , .Q ( coeficiente_b11_L_v_out[8] ) , .IN1 ( n1887 ) , .IN3 ( n1885 ) ) ;
AO22X1 U1250 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[7][8] ) , .Q ( n1886 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[6][8] ) ) ;
AO22X1 U1249 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( \pos_L_reg/bank_registro_registros[4][8] ) , .Q ( n1887 ) 
    , .IN4 ( \pos_L_reg/bank_registro_registros[5][8] ) ) ;
OR4X1 U1248 (.IN4 ( n1880 ) , .IN2 ( n1882 ) 
    , .Q ( coeficiente_b11_L_v_out[7] ) , .IN1 ( n1883 ) , .IN3 ( n1881 ) ) ;
OR4X1 U1263 (.IN4 ( n1900 ) , .IN2 ( n1902 ) , .Q ( in_reg_salida_v[11] ) 
    , .IN1 ( n1903 ) , .IN3 ( n1901 ) ) ;
AO22X1 U1262 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( bank_registro_registros[135] ) , .Q ( n1902 ) 
    , .IN4 ( bank_registro_registros[117] ) ) ;
AO22X1 U1261 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( bank_registro_registros[81] ) , .Q ( n1903 ) 
    , .IN4 ( bank_registro_registros[99] ) ) ;
OR4X1 U1260 (.IN4 ( n1896 ) , .IN2 ( n1898 ) , .Q ( in_reg_salida_v[10] ) 
    , .IN1 ( n1899 ) , .IN3 ( n1897 ) ) ;
AO22X1 U1259 (.IN1 ( n2026 ) , .IN3 ( n2025 ) 
    , .IN2 ( bank_registro_registros[134] ) , .Q ( n1898 ) 
    , .IN4 ( bank_registro_registros[116] ) ) ;
AO22X1 U1258 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( bank_registro_registros[80] ) , .Q ( n1899 ) 
    , .IN4 ( bank_registro_registros[98] ) ) ;
OR4X1 U1257 (.IN4 ( n1892 ) , .IN2 ( n1894 ) , .Q ( in_reg_salida_v[0] ) 
    , .IN1 ( n1895 ) , .IN3 ( n1893 ) ) ;
AO22X1 U1256 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( bank_registro_registros[124] ) , .Q ( n1894 ) 
    , .IN4 ( bank_registro_registros[106] ) ) ;
AO22X1 U1271 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( bank_registro_registros[138] ) , .Q ( n1914 ) 
    , .IN4 ( bank_registro_registros[120] ) ) ;
AO22X1 U1270 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( bank_registro_registros[84] ) , .Q ( n1915 ) 
    , .IN4 ( bank_registro_registros[102] ) ) ;
OR4X1 U1269 (.IN4 ( n1908 ) , .IN2 ( n1910 ) , .Q ( in_reg_salida_v[13] ) 
    , .IN1 ( n1911 ) , .IN3 ( n1909 ) ) ;
AO22X1 U1268 (.IN1 ( n2026 ) , .IN3 ( n2025 ) 
    , .IN2 ( bank_registro_registros[137] ) , .Q ( n1910 ) 
    , .IN4 ( bank_registro_registros[119] ) ) ;
AO22X1 U1267 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( bank_registro_registros[83] ) , .Q ( n1911 ) 
    , .IN4 ( bank_registro_registros[101] ) ) ;
OR4X1 U1266 (.IN4 ( n1904 ) , .IN2 ( n1906 ) , .Q ( in_reg_salida_v[12] ) 
    , .IN1 ( n1907 ) , .IN3 ( n1905 ) ) ;
AO22X1 U1265 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( bank_registro_registros[136] ) , .Q ( n1906 ) 
    , .IN4 ( bank_registro_registros[118] ) ) ;
AO22X1 U1264 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( bank_registro_registros[82] ) , .Q ( n1907 ) 
    , .IN4 ( bank_registro_registros[100] ) ) ;
AO22X1 U1279 (.IN1 ( n1630 ) , .IN3 ( n1633 ) 
    , .IN2 ( bank_registro_registros[123] ) , .Q ( n1927 ) 
    , .IN4 ( bank_registro_registros[33] ) ) ;
NAND4X0 U1278 (.IN1 ( n1925 ) , .QN ( in_reg_salida_v[16] ) , .IN2 ( n1924 ) 
    , .IN3 ( n1931 ) , .IN4 ( n1923 ) ) ;
NOR2X0 U1277 (.QN ( n1924 ) , .IN1 ( n1922 ) , .IN2 ( n1921 ) ) ;
AO22X1 U1276 (.IN1 ( n1630 ) , .IN3 ( n2027 ) 
    , .IN2 ( bank_registro_registros[122] ) , .Q ( n1922 ) 
    , .IN4 ( bank_registro_registros[32] ) ) ;
NAND4X0 U1275 (.IN1 ( n1920 ) , .QN ( in_reg_salida_v[15] ) , .IN2 ( n1919 ) 
    , .IN3 ( n1931 ) , .IN4 ( n1918 ) ) ;
NOR2X0 U1274 (.QN ( n1919 ) , .IN1 ( n1917 ) , .IN2 ( n1916 ) ) ;
AO22X1 U1273 (.IN1 ( n1630 ) , .IN3 ( n2027 ) 
    , .IN2 ( bank_registro_registros[121] ) , .Q ( n1917 ) 
    , .IN4 ( bank_registro_registros[31] ) ) ;
OR4X1 U1272 (.IN4 ( n1912 ) , .IN2 ( n1914 ) , .Q ( in_reg_salida_v[14] ) 
    , .IN1 ( n1915 ) , .IN3 ( n1913 ) ) ;
OR4X1 U1287 (.IN4 ( n1936 ) , .IN2 ( n1938 ) , .Q ( in_reg_salida_v[2] ) 
    , .IN1 ( n1939 ) , .IN3 ( n1937 ) ) ;
AO22X1 U1286 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( bank_registro_registros[126] ) , .Q ( n1938 ) 
    , .IN4 ( bank_registro_registros[108] ) ) ;
AO22X1 U1285 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( bank_registro_registros[72] ) , .Q ( n1939 ) 
    , .IN4 ( bank_registro_registros[90] ) ) ;
OR4X1 U1284 (.IN4 ( n1932 ) , .IN2 ( n1934 ) , .Q ( in_reg_salida_v[1] ) 
    , .IN1 ( n1935 ) , .IN3 ( n1933 ) ) ;
AO22X1 U1283 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( bank_registro_registros[125] ) , .Q ( n1934 ) 
    , .IN4 ( bank_registro_registros[107] ) ) ;
AO22X1 U1282 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( bank_registro_registros[71] ) , .Q ( n1935 ) 
    , .IN4 ( bank_registro_registros[89] ) ) ;
NAND4X0 U1281 (.IN1 ( n1930 ) , .QN ( in_reg_salida_v[17] ) , .IN2 ( n1929 ) 
    , .IN3 ( n1931 ) , .IN4 ( n1928 ) ) ;
NOR2X0 U1280 (.QN ( n1929 ) , .IN1 ( n1927 ) , .IN2 ( n1926 ) ) ;
AO22X1 U1295 (.IN1 ( n1636 ) , .IN3 ( n2027 ) 
    , .IN2 ( bank_registro_registros[5] ) , .Q ( n1949 ) 
    , .IN4 ( bank_registro_registros[21] ) ) ;
AO22X1 U1294 (.IN1 ( n1631 ) , .IN3 ( n2025 ) 
    , .IN2 ( bank_registro_registros[129] ) , .Q ( n1950 ) 
    , .IN4 ( bank_registro_registros[111] ) ) ;
OR4X1 U1293 (.IN4 ( n1944 ) , .IN2 ( n1946 ) , .Q ( in_reg_salida_v[4] ) 
    , .IN1 ( n1947 ) , .IN3 ( n1945 ) ) ;
AO22X1 U1292 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( bank_registro_registros[128] ) , .Q ( n1946 ) 
    , .IN4 ( bank_registro_registros[110] ) ) ;
AO22X1 U1291 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( bank_registro_registros[74] ) , .Q ( n1947 ) 
    , .IN4 ( bank_registro_registros[92] ) ) ;
OR4X1 U1290 (.IN4 ( n1940 ) , .IN2 ( n1942 ) , .Q ( in_reg_salida_v[3] ) 
    , .IN1 ( n1943 ) , .IN3 ( n1941 ) ) ;
AO22X1 U1289 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( bank_registro_registros[127] ) , .Q ( n1942 ) 
    , .IN4 ( bank_registro_registros[109] ) ) ;
AO22X1 U1288 (.IN1 ( n1628 ) , .IN3 ( n1627 ) 
    , .IN2 ( bank_registro_registros[73] ) , .Q ( n1943 ) 
    , .IN4 ( bank_registro_registros[91] ) ) ;
AO22X1 U1303 (.IN1 ( n1631 ) , .IN3 ( n2025 ) 
    , .IN2 ( bank_registro_registros[132] ) , .Q ( n1962 ) 
    , .IN4 ( bank_registro_registros[114] ) ) ;
OR4X1 U1302 (.IN4 ( n1956 ) , .IN2 ( n1958 ) , .Q ( in_reg_salida_v[7] ) 
    , .IN1 ( n1959 ) , .IN3 ( n1957 ) ) ;
AO22X1 U1301 (.IN1 ( n1636 ) , .IN3 ( n2027 ) 
    , .IN2 ( bank_registro_registros[7] ) , .Q ( n1957 ) 
    , .IN4 ( bank_registro_registros[23] ) ) ;
AO22X1 U1300 (.IN1 ( n1631 ) , .IN3 ( n2025 ) 
    , .IN2 ( bank_registro_registros[131] ) , .Q ( n1958 ) 
    , .IN4 ( bank_registro_registros[113] ) ) ;
OR4X1 U1299 (.IN4 ( n1952 ) , .IN2 ( n1954 ) , .Q ( in_reg_salida_v[6] ) 
    , .IN1 ( n1955 ) , .IN3 ( n1953 ) ) ;
AO22X1 U1298 (.IN1 ( n1636 ) , .IN3 ( n2027 ) 
    , .IN2 ( bank_registro_registros[6] ) , .Q ( n1953 ) 
    , .IN4 ( bank_registro_registros[22] ) ) ;
AO22X1 U1297 (.IN1 ( n2026 ) , .IN3 ( n1629 ) 
    , .IN2 ( bank_registro_registros[130] ) , .Q ( n1954 ) 
    , .IN4 ( bank_registro_registros[112] ) ) ;
OR4X1 U1296 (.IN4 ( n1948 ) , .IN2 ( n1950 ) , .Q ( in_reg_salida_v[5] ) 
    , .IN1 ( n1951 ) , .IN3 ( n1949 ) ) ;
AO22X1 U1311 (.IN1 ( n1631 ) , .IN3 ( n1629 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[7][11] ) , .Q ( n1974 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[6][11] ) ) ;
AO22X1 U1310 (.IN1 ( n1636 ) , .IN3 ( n2027 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[0][10] ) , .Q ( n1969 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[1][10] ) ) ;
AO22X1 U1309 (.IN1 ( n1631 ) , .IN3 ( n2025 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[7][10] ) , .Q ( n1970 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[6][10] ) ) ;
OR4X1 U1308 (.IN4 ( n1964 ) , .IN2 ( n1966 ) , .Q ( in_reg_salida_v[9] ) 
    , .IN1 ( n1967 ) , .IN3 ( n1965 ) ) ;
AO22X1 U1307 (.IN1 ( n1636 ) , .IN3 ( n2027 ) 
    , .IN2 ( bank_registro_registros[9] ) , .Q ( n1965 ) 
    , .IN4 ( bank_registro_registros[25] ) ) ;
AO22X1 U1306 (.IN1 ( n1631 ) , .IN3 ( n2025 ) 
    , .IN2 ( bank_registro_registros[133] ) , .Q ( n1966 ) 
    , .IN4 ( bank_registro_registros[115] ) ) ;
OR4X1 U1305 (.IN4 ( n1960 ) , .IN2 ( n1962 ) , .Q ( in_reg_salida_v[8] ) 
    , .IN1 ( n1963 ) , .IN3 ( n1961 ) ) ;
AO22X1 U1304 (.IN1 ( n1636 ) , .IN3 ( n2027 ) 
    , .IN2 ( bank_registro_registros[8] ) , .Q ( n1961 ) 
    , .IN4 ( bank_registro_registros[24] ) ) ;
AO22X1 U1319 (.IN1 ( n1631 ) , .IN3 ( n1629 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[7][15] ) , .Q ( n1990 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[6][15] ) ) ;
AO22X1 U1318 (.IN1 ( n1636 ) , .IN3 ( n1633 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[0][14] ) , .Q ( n1985 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[1][14] ) ) ;
AO22X1 U1317 (.IN1 ( n1631 ) , .IN3 ( n1629 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[7][14] ) , .Q ( n1986 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[6][14] ) ) ;
AO22X1 U1316 (.IN1 ( n1636 ) , .IN3 ( n2027 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[0][13] ) , .Q ( n1981 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[1][13] ) ) ;
AO22X1 U1315 (.IN1 ( n1631 ) , .IN3 ( n2025 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[7][13] ) , .Q ( n1982 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[6][13] ) ) ;
AO22X1 U1314 (.IN1 ( n1636 ) , .IN3 ( n2027 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[0][12] ) , .Q ( n1977 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[1][12] ) ) ;
AO22X1 U1313 (.IN1 ( n1631 ) , .IN3 ( n1629 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[7][12] ) , .Q ( n1978 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[6][12] ) ) ;
AO22X1 U1312 (.IN1 ( n1636 ) , .IN3 ( n2027 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[0][11] ) , .Q ( n1973 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[1][11] ) ) ;
AO22X1 U1327 (.IN1 ( n1636 ) , .IN3 ( n1633 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[0][5] ) , .Q ( n2009 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[1][5] ) ) ;
AO22X1 U1326 (.IN1 ( n2026 ) , .IN3 ( n1629 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[7][5] ) , .Q ( n2010 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[6][5] ) ) ;
AO22X1 U1325 (.IN1 ( n1636 ) , .IN3 ( n1633 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[0][4] ) , .Q ( n2005 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[1][4] ) ) ;
AO22X1 U1324 (.IN1 ( n2026 ) , .IN3 ( n1629 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[7][4] ) , .Q ( n2006 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[6][4] ) ) ;
AO22X1 U1323 (.IN1 ( n1631 ) , .IN3 ( n1629 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[7][18] ) , .Q ( n2002 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[6][18] ) ) ;
AO22X1 U1322 (.IN1 ( n1631 ) , .IN3 ( n1629 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[7][17] ) , .Q ( n1998 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[6][17] ) ) ;
AO22X1 U1321 (.IN1 ( n1631 ) , .IN3 ( n1629 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[7][16] ) , .Q ( n1994 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[6][16] ) ) ;
AO22X1 U1320 (.IN1 ( n1636 ) , .IN3 ( n1633 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[0][15] ) , .Q ( n1989 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[1][15] ) ) ;
AO22X1 U1335 (.IN1 ( n1632 ) , .IN3 ( n2025 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[7][9] ) , .Q ( n2033 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[6][9] ) ) ;
AO22X1 U1334 (.IN1 ( n1628 ) , .IN3 ( n1626 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[4][9] ) , .Q ( n2034 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[5][9] ) ) ;
AO22X1 U1333 (.IN1 ( n1636 ) , .IN3 ( n1633 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[0][8] ) , .Q ( n2021 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[1][8] ) ) ;
AO22X1 U1332 (.IN1 ( n1631 ) , .IN3 ( n1629 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[7][8] ) , .Q ( n2022 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[6][8] ) ) ;
AO22X1 U1331 (.IN1 ( n1636 ) , .IN3 ( n1633 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[0][7] ) , .Q ( n2017 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[1][7] ) ) ;
AO22X1 U1330 (.IN1 ( n1631 ) , .IN3 ( n1629 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[7][7] ) , .Q ( n2018 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[6][7] ) ) ;
AO22X1 U1329 (.IN1 ( n1636 ) , .IN3 ( n1633 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[0][6] ) , .Q ( n2013 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[1][6] ) ) ;
AO22X1 U1328 (.IN1 ( n2026 ) , .IN3 ( n1629 ) 
    , .IN2 ( \sos1_reg/bank_registro_registros[7][6] ) , .Q ( n2014 ) 
    , .IN4 ( \sos1_reg/bank_registro_registros[6][6] ) ) ;
endmodule
